##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Wed Dec 15 22:19:56 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERctr
  CLASS BLOCK ;
  SIZE 70.800000 BY 40.800000 ;
  FOREIGN BATCHARGERctr 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN cc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.720000 40.160000 1.880000 40.800000 ;
    END
  END cc
  PIN tc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 27.320000 40.160000 27.480000 40.800000 ;
    END
  END tc
  PIN cv
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.320000 40.160000 3.480000 40.800000 ;
    END
  END cv
  PIN imonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 19.320000 40.160000 19.480000 40.800000 ;
    END
  END imonen
  PIN vmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 60.920000 40.160000 61.080000 40.800000 ;
    END
  END vmonen
  PIN tmonen
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 47.320000 40.160000 47.480000 40.800000 ;
    END
  END tmonen
  PIN vtok
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 68.120000 40.160000 68.280000 40.800000 ;
    END
  END vtok
  PIN vbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 53.720000 40.160000 53.880000 40.800000 ;
    END
  END vbat[7]
  PIN vbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 52.920000 40.160000 53.080000 40.800000 ;
    END
  END vbat[6]
  PIN vbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 52.120000 40.160000 52.280000 40.800000 ;
    END
  END vbat[5]
  PIN vbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 51.320000 40.160000 51.480000 40.800000 ;
    END
  END vbat[4]
  PIN vbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 50.520000 40.160000 50.680000 40.800000 ;
    END
  END vbat[3]
  PIN vbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 49.720000 40.160000 49.880000 40.800000 ;
    END
  END vbat[2]
  PIN vbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.920000 40.160000 49.080000 40.800000 ;
    END
  END vbat[1]
  PIN vbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 48.120000 40.160000 48.280000 40.800000 ;
    END
  END vbat[0]
  PIN ibat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.120000 40.160000 12.280000 40.800000 ;
    END
  END ibat[7]
  PIN ibat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 11.320000 40.160000 11.480000 40.800000 ;
    END
  END ibat[6]
  PIN ibat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.520000 40.160000 10.680000 40.800000 ;
    END
  END ibat[5]
  PIN ibat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.720000 40.160000 9.880000 40.800000 ;
    END
  END ibat[4]
  PIN ibat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 8.920000 40.160000 9.080000 40.800000 ;
    END
  END ibat[3]
  PIN ibat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 8.120000 40.160000 8.280000 40.800000 ;
    END
  END ibat[2]
  PIN ibat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.320000 40.160000 7.480000 40.800000 ;
    END
  END ibat[1]
  PIN ibat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.520000 40.160000 6.680000 40.800000 ;
    END
  END ibat[0]
  PIN tbat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 26.520000 40.160000 26.680000 40.800000 ;
    END
  END tbat[7]
  PIN tbat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 25.720000 40.160000 25.880000 40.800000 ;
    END
  END tbat[6]
  PIN tbat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.920000 40.160000 25.080000 40.800000 ;
    END
  END tbat[5]
  PIN tbat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.120000 40.160000 24.280000 40.800000 ;
    END
  END tbat[4]
  PIN tbat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 23.320000 40.160000 23.480000 40.800000 ;
    END
  END tbat[3]
  PIN tbat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 22.520000 40.160000 22.680000 40.800000 ;
    END
  END tbat[2]
  PIN tbat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 21.720000 40.160000 21.880000 40.800000 ;
    END
  END tbat[1]
  PIN tbat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 20.920000 40.160000 21.080000 40.800000 ;
    END
  END tbat[0]
  PIN vcutoff[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 60.120000 40.160000 60.280000 40.800000 ;
    END
  END vcutoff[7]
  PIN vcutoff[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 59.320000 40.160000 59.480000 40.800000 ;
    END
  END vcutoff[6]
  PIN vcutoff[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 58.520000 40.160000 58.680000 40.800000 ;
    END
  END vcutoff[5]
  PIN vcutoff[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 57.720000 40.160000 57.880000 40.800000 ;
    END
  END vcutoff[4]
  PIN vcutoff[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 56.920000 40.160000 57.080000 40.800000 ;
    END
  END vcutoff[3]
  PIN vcutoff[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 56.120000 40.160000 56.280000 40.800000 ;
    END
  END vcutoff[2]
  PIN vcutoff[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 55.320000 40.160000 55.480000 40.800000 ;
    END
  END vcutoff[1]
  PIN vcutoff[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 54.520000 40.160000 54.680000 40.800000 ;
    END
  END vcutoff[0]
  PIN vpreset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 67.320000 40.160000 67.480000 40.800000 ;
    END
  END vpreset[7]
  PIN vpreset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 66.520000 40.160000 66.680000 40.800000 ;
    END
  END vpreset[6]
  PIN vpreset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 65.720000 40.160000 65.880000 40.800000 ;
    END
  END vpreset[5]
  PIN vpreset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 64.920000 40.160000 65.080000 40.800000 ;
    END
  END vpreset[4]
  PIN vpreset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 64.120000 40.160000 64.280000 40.800000 ;
    END
  END vpreset[3]
  PIN vpreset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.320000 40.160000 63.480000 40.800000 ;
    END
  END vpreset[2]
  PIN vpreset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 62.520000 40.160000 62.680000 40.800000 ;
    END
  END vpreset[1]
  PIN vpreset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 61.720000 40.160000 61.880000 40.800000 ;
    END
  END vpreset[0]
  PIN tempmin[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 40.120000 40.160000 40.280000 40.800000 ;
    END
  END tempmin[7]
  PIN tempmin[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 39.320000 40.160000 39.480000 40.800000 ;
    END
  END tempmin[6]
  PIN tempmin[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 38.520000 40.160000 38.680000 40.800000 ;
    END
  END tempmin[5]
  PIN tempmin[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 37.720000 40.160000 37.880000 40.800000 ;
    END
  END tempmin[4]
  PIN tempmin[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 36.920000 40.160000 37.080000 40.800000 ;
    END
  END tempmin[3]
  PIN tempmin[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 36.120000 40.160000 36.280000 40.800000 ;
    END
  END tempmin[2]
  PIN tempmin[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 35.320000 40.160000 35.480000 40.800000 ;
    END
  END tempmin[1]
  PIN tempmin[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 34.520000 40.160000 34.680000 40.800000 ;
    END
  END tempmin[0]
  PIN tempmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 33.720000 40.160000 33.880000 40.800000 ;
    END
  END tempmax[7]
  PIN tempmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 32.920000 40.160000 33.080000 40.800000 ;
    END
  END tempmax[6]
  PIN tempmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 32.120000 40.160000 32.280000 40.800000 ;
    END
  END tempmax[5]
  PIN tempmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 31.320000 40.160000 31.480000 40.800000 ;
    END
  END tempmax[4]
  PIN tempmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.520000 40.160000 30.680000 40.800000 ;
    END
  END tempmax[3]
  PIN tempmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 29.720000 40.160000 29.880000 40.800000 ;
    END
  END tempmax[2]
  PIN tempmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.920000 40.160000 29.080000 40.800000 ;
    END
  END tempmax[1]
  PIN tempmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.120000 40.160000 28.280000 40.800000 ;
    END
  END tempmax[0]
  PIN tmax[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 46.520000 40.160000 46.680000 40.800000 ;
    END
  END tmax[7]
  PIN tmax[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 45.720000 40.160000 45.880000 40.800000 ;
    END
  END tmax[6]
  PIN tmax[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 44.920000 40.160000 45.080000 40.800000 ;
    END
  END tmax[5]
  PIN tmax[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 44.120000 40.160000 44.280000 40.800000 ;
    END
  END tmax[4]
  PIN tmax[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 43.320000 40.160000 43.480000 40.800000 ;
    END
  END tmax[3]
  PIN tmax[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 42.520000 40.160000 42.680000 40.800000 ;
    END
  END tmax[2]
  PIN tmax[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 41.720000 40.160000 41.880000 40.800000 ;
    END
  END tmax[1]
  PIN tmax[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 40.920000 40.160000 41.080000 40.800000 ;
    END
  END tmax[0]
  PIN iend[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.520000 40.160000 18.680000 40.800000 ;
    END
  END iend[7]
  PIN iend[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 17.720000 40.160000 17.880000 40.800000 ;
    END
  END iend[6]
  PIN iend[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 16.920000 40.160000 17.080000 40.800000 ;
    END
  END iend[5]
  PIN iend[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 16.120000 40.160000 16.280000 40.800000 ;
    END
  END iend[4]
  PIN iend[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.320000 40.160000 15.480000 40.800000 ;
    END
  END iend[3]
  PIN iend[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 14.520000 40.160000 14.680000 40.800000 ;
    END
  END iend[2]
  PIN iend[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 13.720000 40.160000 13.880000 40.800000 ;
    END
  END iend[1]
  PIN iend[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.920000 40.160000 13.080000 40.800000 ;
    END
  END iend[0]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.520000 40.160000 2.680000 40.800000 ;
    END
  END clk
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.720000 40.160000 5.880000 40.800000 ;
    END
  END en
  PIN rstz
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 20.120000 40.160000 20.280000 40.800000 ;
    END
  END rstz
  PIN dvdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 20.500000 0.640000 21.500000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 0.100000 0.640000 1.100000 ;
    END
  END dgnd
  OBS
    LAYER metal1 ;
      RECT 68.440000 40.000000 70.800000 40.800000 ;
      RECT 67.640000 40.000000 67.960000 40.800000 ;
      RECT 66.840000 40.000000 67.160000 40.800000 ;
      RECT 66.040000 40.000000 66.360000 40.800000 ;
      RECT 65.240000 40.000000 65.560000 40.800000 ;
      RECT 64.440000 40.000000 64.760000 40.800000 ;
      RECT 63.640000 40.000000 63.960000 40.800000 ;
      RECT 62.840000 40.000000 63.160000 40.800000 ;
      RECT 62.040000 40.000000 62.360000 40.800000 ;
      RECT 61.240000 40.000000 61.560000 40.800000 ;
      RECT 60.440000 40.000000 60.760000 40.800000 ;
      RECT 59.640000 40.000000 59.960000 40.800000 ;
      RECT 58.840000 40.000000 59.160000 40.800000 ;
      RECT 58.040000 40.000000 58.360000 40.800000 ;
      RECT 57.240000 40.000000 57.560000 40.800000 ;
      RECT 56.440000 40.000000 56.760000 40.800000 ;
      RECT 55.640000 40.000000 55.960000 40.800000 ;
      RECT 54.840000 40.000000 55.160000 40.800000 ;
      RECT 54.040000 40.000000 54.360000 40.800000 ;
      RECT 53.240000 40.000000 53.560000 40.800000 ;
      RECT 52.440000 40.000000 52.760000 40.800000 ;
      RECT 51.640000 40.000000 51.960000 40.800000 ;
      RECT 50.840000 40.000000 51.160000 40.800000 ;
      RECT 50.040000 40.000000 50.360000 40.800000 ;
      RECT 49.240000 40.000000 49.560000 40.800000 ;
      RECT 48.440000 40.000000 48.760000 40.800000 ;
      RECT 47.640000 40.000000 47.960000 40.800000 ;
      RECT 46.840000 40.000000 47.160000 40.800000 ;
      RECT 46.040000 40.000000 46.360000 40.800000 ;
      RECT 45.240000 40.000000 45.560000 40.800000 ;
      RECT 44.440000 40.000000 44.760000 40.800000 ;
      RECT 43.640000 40.000000 43.960000 40.800000 ;
      RECT 42.840000 40.000000 43.160000 40.800000 ;
      RECT 42.040000 40.000000 42.360000 40.800000 ;
      RECT 41.240000 40.000000 41.560000 40.800000 ;
      RECT 40.440000 40.000000 40.760000 40.800000 ;
      RECT 39.640000 40.000000 39.960000 40.800000 ;
      RECT 38.840000 40.000000 39.160000 40.800000 ;
      RECT 38.040000 40.000000 38.360000 40.800000 ;
      RECT 37.240000 40.000000 37.560000 40.800000 ;
      RECT 36.440000 40.000000 36.760000 40.800000 ;
      RECT 35.640000 40.000000 35.960000 40.800000 ;
      RECT 34.840000 40.000000 35.160000 40.800000 ;
      RECT 34.040000 40.000000 34.360000 40.800000 ;
      RECT 33.240000 40.000000 33.560000 40.800000 ;
      RECT 32.440000 40.000000 32.760000 40.800000 ;
      RECT 31.640000 40.000000 31.960000 40.800000 ;
      RECT 30.840000 40.000000 31.160000 40.800000 ;
      RECT 30.040000 40.000000 30.360000 40.800000 ;
      RECT 29.240000 40.000000 29.560000 40.800000 ;
      RECT 28.440000 40.000000 28.760000 40.800000 ;
      RECT 27.640000 40.000000 27.960000 40.800000 ;
      RECT 26.840000 40.000000 27.160000 40.800000 ;
      RECT 26.040000 40.000000 26.360000 40.800000 ;
      RECT 25.240000 40.000000 25.560000 40.800000 ;
      RECT 24.440000 40.000000 24.760000 40.800000 ;
      RECT 23.640000 40.000000 23.960000 40.800000 ;
      RECT 22.840000 40.000000 23.160000 40.800000 ;
      RECT 22.040000 40.000000 22.360000 40.800000 ;
      RECT 21.240000 40.000000 21.560000 40.800000 ;
      RECT 20.440000 40.000000 20.760000 40.800000 ;
      RECT 19.640000 40.000000 19.960000 40.800000 ;
      RECT 18.840000 40.000000 19.160000 40.800000 ;
      RECT 18.040000 40.000000 18.360000 40.800000 ;
      RECT 17.240000 40.000000 17.560000 40.800000 ;
      RECT 16.440000 40.000000 16.760000 40.800000 ;
      RECT 15.640000 40.000000 15.960000 40.800000 ;
      RECT 14.840000 40.000000 15.160000 40.800000 ;
      RECT 14.040000 40.000000 14.360000 40.800000 ;
      RECT 13.240000 40.000000 13.560000 40.800000 ;
      RECT 12.440000 40.000000 12.760000 40.800000 ;
      RECT 11.640000 40.000000 11.960000 40.800000 ;
      RECT 10.840000 40.000000 11.160000 40.800000 ;
      RECT 10.040000 40.000000 10.360000 40.800000 ;
      RECT 9.240000 40.000000 9.560000 40.800000 ;
      RECT 8.440000 40.000000 8.760000 40.800000 ;
      RECT 7.640000 40.000000 7.960000 40.800000 ;
      RECT 6.840000 40.000000 7.160000 40.800000 ;
      RECT 6.040000 40.000000 6.360000 40.800000 ;
      RECT 3.640000 40.000000 5.560000 40.800000 ;
      RECT 2.840000 40.000000 3.160000 40.800000 ;
      RECT 2.040000 40.000000 2.360000 40.800000 ;
      RECT 0.000000 40.000000 1.560000 40.800000 ;
      RECT 0.000000 21.660000 70.800000 40.000000 ;
      RECT 0.800000 20.340000 70.800000 21.660000 ;
      RECT 0.000000 1.260000 70.800000 20.340000 ;
      RECT 0.800000 0.000000 70.800000 1.260000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 70.800000 40.800000 ;
  END
END BATCHARGERctr

END LIBRARY
