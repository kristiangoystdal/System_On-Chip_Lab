##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Sun Dec 19 17:29:01 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO FULLCHIPcore
  CLASS BLOCK ;
  SIZE 50.000000 BY 76.800000 ;
  FOREIGN FULLCHIPcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN count_dir
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 42.000000 0.260000 42.400000 ;
    END
  END count_dir
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 46.000000 0.260000 46.400000 ;
    END
  END enable
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 50.000000 0.260000 50.400000 ;
    END
  END reset
  PIN count[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 38.000000 0.260000 38.400000 ;
    END
  END count[3]
  PIN count[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 34.000000 0.260000 34.400000 ;
    END
  END count[2]
  PIN count[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 30.000000 0.260000 30.400000 ;
    END
  END count[1]
  PIN count[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 26.000000 0.260000 26.400000 ;
    END
  END count[0]
  PIN vctrl
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER metal1 ;
        RECT 49.740000 30.000000 50.000000 30.400000 ;
    END
  END vctrl
  PIN avdd
    DIRECTION INOUT ;
#    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 49.840000 53.600000 50.000000 55.600000 ;
    END
  END avdd
  PIN agnd
    DIRECTION INOUT ;
#    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 49.840000 3.200000 50.000000 5.200000 ;
    END
  END agnd
  PIN dvdd
    DIRECTION INOUT ;
#    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 49.840000 20.800000 50.000000 22.800000 ;
    END
  END dvdd
  OBS
    LAYER metal1 ;
      RECT 0.000000 50.560000 50.000000 76.800000 ;
      RECT 0.420000 49.840000 50.000000 50.560000 ;
      RECT 0.000000 46.560000 50.000000 49.840000 ;
      RECT 0.420000 45.840000 50.000000 46.560000 ;
      RECT 0.000000 42.560000 50.000000 45.840000 ;
      RECT 0.420000 41.840000 50.000000 42.560000 ;
      RECT 0.000000 38.560000 50.000000 41.840000 ;
      RECT 0.420000 37.840000 50.000000 38.560000 ;
      RECT 0.000000 34.560000 50.000000 37.840000 ;
      RECT 0.420000 33.840000 50.000000 34.560000 ;
      RECT 0.000000 30.560000 50.000000 33.840000 ;
      RECT 0.420000 29.840000 49.580000 30.560000 ;
      RECT 0.000000 26.560000 50.000000 29.840000 ;
      RECT 0.420000 25.840000 50.000000 26.560000 ;
      RECT 0.000000 0.000000 50.000000 25.840000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 50.000000 76.800000 ;
    LAYER metal3 ;
      RECT 0.000000 55.880000 50.000000 76.800000 ;
      RECT 0.000000 53.320000 49.560000 55.880000 ;
      RECT 0.000000 23.080000 50.000000 53.320000 ;
      RECT 0.000000 20.520000 49.560000 23.080000 ;
      RECT 0.000000 5.480000 50.000000 20.520000 ;
      RECT 0.000000 2.920000 49.560000 5.480000 ;
      RECT 0.000000 0.000000 50.000000 2.920000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 50.000000 76.800000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 50.000000 76.800000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 50.000000 76.800000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 50.000000 76.800000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 50.000000 76.800000 ;
  END
END FULLCHIPcore

END LIBRARY
