##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Wed Dec 15 20:04:39 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERsaradc
  CLASS BLOCK ;
  SIZE 200.800000 BY 120.800000 ;
  FOREIGN BATCHARGERsaradc 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN vbat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 134.520000 0.000000 134.680000 0.640000 ;
    END
  END vbat[7]
  PIN vbat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 138.520000 0.000000 138.680000 0.640000 ;
    END
  END vbat[6]
  PIN vbat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 142.520000 0.000000 142.680000 0.640000 ;
    END
  END vbat[5]
  PIN vbat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 146.520000 0.000000 146.680000 0.640000 ;
    END
  END vbat[4]
  PIN vbat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 150.520000 0.000000 150.680000 0.640000 ;
    END
  END vbat[3]
  PIN vbat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 154.520000 0.000000 154.680000 0.640000 ;
    END
  END vbat[2]
  PIN vbat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 158.520000 0.000000 158.680000 0.640000 ;
    END
  END vbat[1]
  PIN vbat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 162.520000 0.000000 162.680000 0.640000 ;
    END
  END vbat[0]
  PIN ibat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 130.120000 120.160000 130.280000 120.800000 ;
    END
  END ibat[7]
  PIN ibat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 120.120000 120.160000 120.280000 120.800000 ;
    END
  END ibat[6]
  PIN ibat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 110.120000 120.160000 110.280000 120.800000 ;
    END
  END ibat[5]
  PIN ibat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 100.120000 120.160000 100.280000 120.800000 ;
    END
  END ibat[4]
  PIN ibat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 90.120000 120.160000 90.280000 120.800000 ;
    END
  END ibat[3]
  PIN ibat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 80.120000 120.160000 80.280000 120.800000 ;
    END
  END ibat[2]
  PIN ibat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 70.120000 120.160000 70.280000 120.800000 ;
    END
  END ibat[1]
  PIN ibat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 60.120000 120.160000 60.280000 120.800000 ;
    END
  END ibat[0]
  PIN tbat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 170.520000 0.000000 170.680000 0.640000 ;
    END
  END tbat[7]
  PIN tbat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 174.520000 0.000000 174.680000 0.640000 ;
    END
  END tbat[6]
  PIN tbat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 178.520000 0.000000 178.680000 0.640000 ;
    END
  END tbat[5]
  PIN tbat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 182.520000 0.000000 182.680000 0.640000 ;
    END
  END tbat[4]
  PIN tbat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 186.520000 0.000000 186.680000 0.640000 ;
    END
  END tbat[3]
  PIN tbat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 190.520000 0.000000 190.680000 0.640000 ;
    END
  END tbat[2]
  PIN tbat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 194.520000 0.000000 194.680000 0.640000 ;
    END
  END tbat[1]
  PIN tbat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 198.520000 0.000000 198.680000 0.640000 ;
    END
  END tbat[0]
  PIN vtok
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 110.520000 0.000000 110.680000 0.640000 ;
    END
  END vtok
  PIN vref
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 114.520000 0.000000 114.680000 0.640000 ;
    END
  END vref
  PIN ibias1u
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 140.120000 120.160000 140.280000 120.800000 ;
    END
  END ibias1u
  PIN vbattemp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 126.520000 0.000000 126.680000 0.640000 ;
    END
  END vbattemp
  PIN vbatvolt
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 122.520000 0.000000 122.680000 0.640000 ;
    END
  END vbatvolt
  PIN vbatcurr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 130.520000 0.000000 130.680000 0.640000 ;
    END
  END vbatcurr
  PIN imeasen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 150.120000 120.160000 150.280000 120.800000 ;
    END
  END imeasen
  PIN vmeasen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 118.520000 0.000000 118.680000 0.640000 ;
    END
  END vmeasen
  PIN tmeasen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 166.520000 0.000000 166.680000 0.640000 ;
    END
  END tmeasen
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 50.120000 120.160000 50.280000 120.800000 ;
    END
  END en
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 72.520000 0.000000 72.680000 0.640000 ;
    END
  END clk
  PIN rstz
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 160.120000 120.160000 160.280000 120.800000 ;
    END
  END rstz
  PIN avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.700000 120.160000 4.700000 120.800000 ;
    END
  END avdd
  PIN dvdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 28.500000 0.000000 29.500000 0.640000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 29.700000 120.160000 30.700000 120.800000 ;
    END
  END dgnd
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.700000 0.000000 2.700000 0.640000 ;
    END
  END agnd
  OBS
    LAYER metal1 ;
      RECT 160.440000 120.000000 200.800000 120.800000 ;
      RECT 150.440000 120.000000 159.960000 120.800000 ;
      RECT 140.440000 120.000000 149.960000 120.800000 ;
      RECT 130.440000 120.000000 139.960000 120.800000 ;
      RECT 120.440000 120.000000 129.960000 120.800000 ;
      RECT 110.440000 120.000000 119.960000 120.800000 ;
      RECT 100.440000 120.000000 109.960000 120.800000 ;
      RECT 90.440000 120.000000 99.960000 120.800000 ;
      RECT 80.440000 120.000000 89.960000 120.800000 ;
      RECT 70.440000 120.000000 79.960000 120.800000 ;
      RECT 60.440000 120.000000 69.960000 120.800000 ;
      RECT 50.440000 120.000000 59.960000 120.800000 ;
      RECT 30.860000 120.000000 49.960000 120.800000 ;
      RECT 4.860000 120.000000 29.540000 120.800000 ;
      RECT 0.000000 120.000000 3.540000 120.800000 ;
      RECT 0.000000 0.800000 200.800000 120.000000 ;
      RECT 198.840000 0.000000 200.800000 0.800000 ;
      RECT 194.840000 0.000000 198.360000 0.800000 ;
      RECT 190.840000 0.000000 194.360000 0.800000 ;
      RECT 186.840000 0.000000 190.360000 0.800000 ;
      RECT 182.840000 0.000000 186.360000 0.800000 ;
      RECT 178.840000 0.000000 182.360000 0.800000 ;
      RECT 174.840000 0.000000 178.360000 0.800000 ;
      RECT 170.840000 0.000000 174.360000 0.800000 ;
      RECT 166.840000 0.000000 170.360000 0.800000 ;
      RECT 162.840000 0.000000 166.360000 0.800000 ;
      RECT 158.840000 0.000000 162.360000 0.800000 ;
      RECT 154.840000 0.000000 158.360000 0.800000 ;
      RECT 150.840000 0.000000 154.360000 0.800000 ;
      RECT 146.840000 0.000000 150.360000 0.800000 ;
      RECT 142.840000 0.000000 146.360000 0.800000 ;
      RECT 138.840000 0.000000 142.360000 0.800000 ;
      RECT 134.840000 0.000000 138.360000 0.800000 ;
      RECT 130.840000 0.000000 134.360000 0.800000 ;
      RECT 126.840000 0.000000 130.360000 0.800000 ;
      RECT 122.840000 0.000000 126.360000 0.800000 ;
      RECT 118.840000 0.000000 122.360000 0.800000 ;
      RECT 114.840000 0.000000 118.360000 0.800000 ;
      RECT 110.840000 0.000000 114.360000 0.800000 ;
      RECT 72.840000 0.000000 110.360000 0.800000 ;
      RECT 29.660000 0.000000 72.360000 0.800000 ;
      RECT 2.860000 0.000000 28.340000 0.800000 ;
      RECT 0.000000 0.000000 1.540000 0.800000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 200.800000 120.800000 ;
  END
END BATCHARGERsaradc

END LIBRARY
