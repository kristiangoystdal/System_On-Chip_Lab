##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Tue Jan  7 12:35:30 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO counter4bit
  CLASS BLOCK ;
  SIZE 29.200000 BY 26.400000 ;
  FOREIGN counter4bit 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 14.900000 0.000000 15.100000 0.520000 ;
    END
  END clk
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 12.900000 0.520000 13.100000 ;
    END
  END enable
  PIN count_dir
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 12.500000 0.520000 12.700000 ;
    END
  END count_dir
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.000000 13.300000 0.520000 13.500000 ;
    END
  END reset
  PIN count[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 28.680000 12.900000 29.200000 13.100000 ;
    END
  END count[3]
  PIN count[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 28.680000 13.300000 29.200000 13.500000 ;
    END
  END count[2]
  PIN count[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 28.680000 13.700000 29.200000 13.900000 ;
    END
  END count[1]
  PIN count[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 28.680000 14.100000 29.200000 14.300000 ;
    END
  END count[0]
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 29.200000 26.400000 ;
    LAYER metal2 ;
      RECT 0.000000 0.720000 29.200000 26.400000 ;
      RECT 15.300000 0.000000 29.200000 0.720000 ;
      RECT 0.000000 0.000000 14.700000 0.720000 ;
    LAYER metal3 ;
      RECT 0.000000 14.500000 29.200000 26.400000 ;
      RECT 0.000000 13.700000 28.480000 14.500000 ;
      RECT 0.720000 12.700000 28.480000 13.700000 ;
      RECT 0.720000 12.300000 29.200000 12.700000 ;
      RECT 0.000000 0.000000 29.200000 12.300000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 29.200000 26.400000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 29.200000 26.400000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 29.200000 26.400000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 29.200000 26.400000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 29.200000 26.400000 ;
  END
END counter4bit

END LIBRARY
