VERSION 5.5 ;
NAMESCASESENSITIVE ON ;

#------------------------------------------
# Preview export LEF
#
#        Preview sub-version 4.4.3.72
#
# TECH LIB NAME: FSC0L_D
# TECH FILE NAME: techfile.cds
# PROCESS OPTION: 8M2T
# DATE : 2004 10 26
#------------------------------------------
 
#------------------------------------------
# case sensitive
#------------------------------------------
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
#------------------------------------------
# declaration of resolution
#------------------------------------------
UNITS
    DATABASE MICRONS 1000  ;
END UNITS
 
MANUFACTURINGGRID 0.01 ;

#------------------------------------------
# declaration of overlap
#------------------------------------------
LAYER overlap
    TYPE OVERLAP ;
END overlap

#------------------------------------------
# declaration of via array spacing 
#------------------------------------------
PROPERTYDEFINITIONS
  LAYER LEF57_SPACING STRING ;
  LAYER LEF57_ARRAYSPACING STRING ;
END PROPERTYDEFINITIONS

#------------------------------------------
# declaration of non-routing layer
#------------------------------------------
#LAYER contact
#    TYPE CUT ;
#END contact

# declaration of routing layer
LAYER metal1
    TYPE ROUTING ;
    WIDTH 0.160 ;
    SPACING 0.160 ;
    SPACING 0.26 RANGE 1.76 1000 ;
    PROPERTY LEF57_SPACING
    "SPACING 0.19 ENDOFLINE 0.181 WITHIN 0.1 PARALLELEDGE 0.19 WITHIN 0.1 TWOEDGES ;" ;
    PITCH 0.400 ;
    OFFSET 0.20 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25 ;
    AREA 0.1024 ;
    MINENCLOSEDAREA 0.3072 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.001047 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    THICKNESS 0.29 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.16 0.32 0.64 1.28 25 ;
    TABLEENTRIES
    21.48 15.82 12.02 9.57 6.45 ;
END metal1

LAYER via
    TYPE CUT ;
    SPACING 0.2 ;
    SPACING 0.28 ADJACENTCUTS 4 WITHIN 0.3 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.28 ARRAYCUTS 3 SPACING 1.2 ;" ;
END via

LAYER metal2
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.200 ;
    SPACING 0.28 RANGE 2 1000 ;
    PITCH 0.400 ;
    OFFSET 0.20 ;
##    WIREEXTENSION 0.16 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25 ;
    AREA 0.1024 ;
    MINENCLOSEDAREA 0.3072 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000913 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    THICKNESS 0.32 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.20 0.40 0.80 1.60 25 ;
    TABLEENTRIES
    13.45 9.64 7.00 5.20 2.54 ;
END metal2

LAYER via2
    TYPE CUT ;
    SPACING 0.2 ;
    SPACING 0.28 ADJACENTCUTS 4 WITHIN 0.3 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.28 ARRAYCUTS 3 SPACING 1.2 ;" ;
END via2

LAYER metal3
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.200 ;
    SPACING 0.28 RANGE 2 1000 ;
    PITCH 0.400 ;
    OFFSET 0.20 ;
##    WIREEXTENSION 0.16 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25 ;
    AREA 0.1024 ;
    MINENCLOSEDAREA 0.3072 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000912 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    THICKNESS 0.32 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.20 0.40 0.80 1.60 25 ;
    TABLEENTRIES
    13.45 9.64 7.00 5.20 2.54 ;
END metal3

LAYER via3
    TYPE CUT ;
    SPACING 0.2 ;
    SPACING 0.28 ADJACENTCUTS 4 WITHIN 0.3 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.28 ARRAYCUTS 3 SPACING 1.2 ;" ;
END via3

LAYER metal4
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.200 ;
    SPACING 0.28 RANGE 2 1000 ;
    PITCH 0.400 ;
    OFFSET 0.20 ;
##    WIREEXTENSION 0.16 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25 ;
    AREA 0.1024 ;
    MINENCLOSEDAREA 0.3072 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000914 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    THICKNESS 0.32 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.20 0.40 0.80 1.60 25 ;
    TABLEENTRIES
    13.45 9.64 7.00 5.20 2.54 ;
END metal4

LAYER via4
    TYPE CUT ;
    SPACING 0.2 ;
    SPACING 0.28 ADJACENTCUTS 4 WITHIN 0.3 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.28 ARRAYCUTS 3 SPACING 1.2 ;" ;
END via4

LAYER metal5
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.200 ;
    SPACING 0.28 RANGE 2 1000 ;
    PITCH 0.400 ;
    OFFSET 0.20 ;
##    WIREEXTENSION 0.16 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25 ;
    AREA 0.1024 ;
    MINENCLOSEDAREA 0.3072 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.000912 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    THICKNESS 0.32 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.20 0.40 0.80 1.60 25 ;
    TABLEENTRIES
    13.45 9.64 7.00 5.20 2.54 ;
END metal5

LAYER via5
    TYPE CUT ;
    SPACING 0.2 ;
    SPACING 0.28 ADJACENTCUTS 4 WITHIN 0.3 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.28 ARRAYCUTS 3 SPACING 1.2 ;" ;
END via5

LAYER metal6
    TYPE ROUTING ;
    WIDTH 0.200 ;
    SPACING 0.200 ;
    SPACING 0.28 RANGE 2 1000 ;
    PITCH 0.400 ;
    OFFSET 0.20 ;
##    WIREEXTENSION 0.16 ;
    MINIMUMCUT 2 WIDTH 1.4 ;
    MAXWIDTH 25 ;
    AREA 0.1024 ;
    MINENCLOSEDAREA 0.3072 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.000914 ;
    RESISTANCE RPERSQ 0.0700000000 ;
    THICKNESS 0.32 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.20 0.40 0.80 1.60 25 ;
    TABLEENTRIES
    13.45 9.64 7.00 5.20 2.54 ;
END metal6

LAYER via6
    TYPE CUT ;
    SPACING 0.4 ;
    SPACING 0.5 ADJACENTCUTS 4 WITHIN 0.7 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.5 ARRAYCUTS 3 SPACING 2.4 ;" ;
END via6
 
LAYER metal7
    TYPE ROUTING ;
    WIDTH 0.400 ;
    SPACING 0.400 ;
    SPACING 0.5 RANGE 1.6 1000 ;
    PITCH 0.800 ;
    OFFSET 0.40 ;
    MAXWIDTH 25 ;
    AREA 0.33 ;
    MINENCLOSEDAREA 0.87 ;
    DIRECTION HORIZONTAL ;
    CAPACITANCE CPERSQDIST 0.00052 ;
    RESISTANCE RPERSQ 0.0270000000 ;
    THICKNESS 0.8 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.40 0.80 1.60 3.20 25 ;
    TABLEENTRIES
    16.90 12.13 8.83 6.59 3.64 ;
END metal7

LAYER via7
    TYPE CUT ;
    SPACING 0.4 ;
    SPACING 0.5 ADJACENTCUTS 4 WITHIN 0.7 ;
    PROPERTY LEF57_ARRAYSPACING
    "ARRAYSPACING WIDTH 5.0 CUTSPACING 0.5 ARRAYCUTS 3 SPACING 2.4 ;" ;
END via7
 
LAYER metal8
    TYPE ROUTING ;
    WIDTH 0.400 ;
    SPACING 0.400 ;
    SPACING 0.5 RANGE 1.6 1000 ;
    PITCH 0.800 ;
    OFFSET 0.40 ;
    MAXWIDTH 25 ;
    AREA 0.33 ;
    MINENCLOSEDAREA 0.87 ;
    DIRECTION VERTICAL ;
    CAPACITANCE CPERSQDIST 0.00047 ;
    RESISTANCE RPERSQ 0.0270000000 ;
    THICKNESS 0.8 ;
    ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH
    0.40 0.80 1.60 3.20 25 ;
    TABLEENTRIES
    16.90 12.13 8.83 6.59 3.64 ;
END metal8

#------------------------------------------
# Define four direction default vias
VIA VIA12_HH DEFAULT
  LAYER metal2 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal1 ;
        RECT -0.16 -0.1 0.16 0.1 ;
END VIA12_HH
VIA VIA12_HV DEFAULT
  LAYER metal2 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal1 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA12_HV
VIA VIA12_VH DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal1 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA12_VH
VIA VIA12_VV DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal1 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA12_VV
VIA VIA23_HH DEFAULT
  LAYER metal2 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA23_HH
VIA VIA23_HV DEFAULT
  LAYER metal2 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA23_HV
VIA VIA23_VH DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA23_VH
VIA VIA23_VV DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA23_VV
VIA VIA34_HH DEFAULT
  LAYER metal4 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA34_HH
VIA VIA34_HV DEFAULT
  LAYER metal4 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA34_HV
VIA VIA34_VH DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA34_VH
VIA VIA34_VV DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal3 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA34_VV
VIA VIA45_HH DEFAULT
  LAYER metal4 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA45_HH
VIA VIA45_HV DEFAULT
  LAYER metal4 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA45_HV
VIA VIA45_VH DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA45_VH
VIA VIA45_VV DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA45_VV
VIA VIA56_HH DEFAULT
  LAYER metal6 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA56_HH
VIA VIA56_HV DEFAULT
  LAYER metal6 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA56_HV
VIA VIA56_VH DEFAULT
  LAYER metal6 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA56_VH
VIA VIA56_VV DEFAULT
  LAYER metal6 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
  LAYER metal5 ;
        RECT -0.1 -0.16 0.1 0.16 ;
  RESISTANCE 1.5 ;
END VIA56_VV
VIA VIA67_Def DEFAULT
  LAYER metal6 ;
        RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via6 ;
        RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
  RESISTANCE 0.6 ;
END VIA67_Def
VIA VIA78_Def DEFAULT
  LAYER metal8 ;
        RECT -0.2 -0.2 0.2 0.2 ;
  LAYER via7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
  LAYER metal7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
  RESISTANCE 0.6 ;
END VIA78_Def
#------------------------------------------


#------------------------------------------
# Define Stack only default vias
VIA VIA23_stack_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER metal2 ;
	 RECT -0.1 -0.36 0.1 0.16 ;
    LAYER via2 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal3 ;
	   RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA23_stack_HAMMER1
VIA VIA23_stack_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER metal2 ;
	 RECT -0.1 -0.16 0.1 0.36 ;
    LAYER via2 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal3 ;
	   RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA23_stack_HAMMER2
VIA VIA23_stack_CROSS DEFAULT TOPOFSTACKONLY
    LAYER metal2 ;
	 RECT -0.1 -0.26 0.1 0.26 ;
    LAYER via2 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal3 ;
	   RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA23_stack_CROSS
VIA VIA34_stack_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER metal4 ;
	   RECT -0.1 -0.16 0.1 0.16 ;
    LAYER via3 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal3 ;
	 RECT -0.36 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA34_stack_HAMMER1
VIA VIA34_stack_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER metal4 ;
	   RECT -0.1 -0.16 0.1 0.16 ;
    LAYER via3 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal3 ;
	 RECT -0.16 -0.1 0.36 0.1 ;
  RESISTANCE 1.5 ;
END VIA34_stack_HAMMER2
VIA VIA34_stack_CROSS DEFAULT TOPOFSTACKONLY
    LAYER metal4 ;
	   RECT -0.1 -0.16 0.1 0.16 ;
    LAYER via3 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal3 ;
	 RECT -0.26 -0.1 0.26 0.1 ;
  RESISTANCE 1.5 ;
END VIA34_stack_CROSS
VIA VIA45_stack_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER metal4 ;
	 RECT -0.1 -0.36 0.1 0.16 ;
    LAYER via4 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal5 ;
	   RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA45_stack_HAMMER1
VIA VIA45_stack_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER metal4 ;
	 RECT -0.1 -0.16 0.1 0.36 ;
    LAYER via4 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal5 ;
	   RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA45_stack_HAMMER2
VIA VIA45_stack_CROSS DEFAULT TOPOFSTACKONLY
    LAYER metal4 ;
	 RECT -0.1 -0.26 0.1 0.26 ;
    LAYER via4 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal5 ;
	   RECT -0.16 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA45_stack_CROSS
VIA VIA56_stack_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER metal6 ;
	   RECT -0.1 -0.16 0.1 0.16 ;
    LAYER via5 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal5 ;
	 RECT -0.36 -0.1 0.16 0.1 ;
  RESISTANCE 1.5 ;
END VIA56_stack_HAMMER1
VIA VIA56_stack_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER metal6 ;
	   RECT -0.1 -0.16 0.1 0.16 ;
    LAYER via5 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal5 ;
	 RECT -0.16 -0.1 0.36 0.1 ;
  RESISTANCE 1.5 ;
END VIA56_stack_HAMMER2
VIA VIA56_stack_CROSS DEFAULT TOPOFSTACKONLY
    LAYER metal6 ;
	   RECT -0.1 -0.16 0.1 0.16 ;
    LAYER via5 ;
	   RECT -0.1 -0.1 0.1 0.1 ;
    LAYER metal5 ;
	 RECT -0.26 -0.1 0.26 0.1 ;
  RESISTANCE 1.5 ;
END VIA56_stack_CROSS
VIA VIA67_stack_Def DEFAULT TOPOFSTACKONLY
    LAYER metal6 ;
	 RECT -0.2 -0.2 0.2 0.2 ;
    LAYER via6 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER metal7 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
  RESISTANCE 0.6 ;
END VIA67_stack_Def
VIA VIA78_stack_HAMMER1 DEFAULT TOPOFSTACKONLY
    LAYER metal8 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER via7 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER metal7 ;
	 RECT -0.63 -0.2 0.2 0.2 ;
  RESISTANCE 0.6 ;
END VIA78_stack_HAMMER1
VIA VIA78_stack_HAMMER2 DEFAULT TOPOFSTACKONLY
    LAYER metal8 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER via7 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER metal7 ;
	 RECT -0.2 -0.2 0.63 0.2 ;
  RESISTANCE 0.6 ;
END VIA78_stack_HAMMER2
VIA VIA78_stack_CROSS DEFAULT TOPOFSTACKONLY
    LAYER metal8 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER via7 ;
	   RECT -0.2 -0.2 0.2 0.2 ;
    LAYER metal7 ;
	 RECT -0.42 -0.2 0.41 0.2 ;
  RESISTANCE 0.6 ;
END VIA78_stack_CROSS
#------------------------------------------

#------------------------------------------
# Define double via for mincut difinition
VIA VIA12_DC_RIGHT DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.5 0.16 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT 0.3 -0.1 0.5 0.1 ;
  LAYER metal1 ;
        RECT -0.16 -0.1 0.56  0.1 ;
END VIA12_DC_RIGHT

VIA VIA12_DC_LEFT DEFAULT
  LAYER metal2 ;
        RECT -0.5 -0.16 0.1 0.16 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.5 -0.1 -0.3 0.1 ;
  LAYER metal1 ;
        RECT -0.56 -0.1 0.16  0.1 ;
END VIA12_DC_LEFT

VIA VIA12_DC_TOP DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.1 0.56 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 0.3 0.1 0.5 ;
  LAYER metal1 ;
        RECT -0.16 -0.1 0.16  0.5 ;
END VIA12_DC_TOP

VIA VIA12_DC_DOWN DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.56 0.1 0.16 ;
  LAYER via ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 -0.5 0.1 -0.3 ;
  LAYER metal1 ;
        RECT -0.16 -0.5 0.16  0.1 ;
END VIA12_DC_DOWN

VIA VIA23_DC_RIGHT DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.5 0.16 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT 0.3 -0.1 0.5 0.1 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.56  0.1 ;
END VIA23_DC_RIGHT

VIA VIA23_DC_LEFT DEFAULT
  LAYER metal2 ;
        RECT -0.5 -0.16 0.1 0.16 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.5 -0.1 -0.3 0.1 ;
  LAYER metal3 ;
        RECT -0.56 -0.1 0.16  0.1 ;
END VIA23_DC_LEFT

VIA VIA23_DC_TOP DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.16 0.1 0.56 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 0.3 0.1 0.5 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.16  0.5 ;
END VIA23_DC_TOP

VIA VIA23_DC_DOWN DEFAULT
  LAYER metal2 ;
        RECT -0.1 -0.56 0.1 0.16 ;
  LAYER via2 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 -0.5 0.1 -0.3 ;
  LAYER metal3 ;
        RECT -0.16 -0.5 0.16  0.1 ;
END VIA23_DC_DOWN

VIA VIA34_DC_RIGHT DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.5 0.16 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT 0.3 -0.1 0.5 0.1 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.56  0.1 ;
END VIA34_DC_RIGHT

VIA VIA34_DC_LEFT DEFAULT
  LAYER metal4 ;
        RECT -0.5 -0.16 0.1 0.16 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.5 -0.1 -0.3 0.1 ;
  LAYER metal3 ;
        RECT -0.56 -0.1 0.16  0.1 ;
END VIA34_DC_LEFT

VIA VIA34_DC_TOP DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.1 0.56 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 0.3 0.1 0.5 ;
  LAYER metal3 ;
        RECT -0.16 -0.1 0.16  0.5 ;
END VIA34_DC_TOP

VIA VIA34_DC_DOWN DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.56 0.1 0.16 ;
  LAYER via3 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 -0.5 0.1 -0.3 ;
  LAYER metal3 ;
        RECT -0.16 -0.5 0.16  0.1 ;
END VIA34_DC_DOWN

VIA VIA45_DC_RIGHT DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.5 0.16 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT 0.3 -0.1 0.5 0.1 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.56  0.1 ;
END VIA45_DC_RIGHT

VIA VIA45_DC_LEFT DEFAULT
  LAYER metal4 ;
        RECT -0.5 -0.16 0.1 0.16 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.5 -0.1 -0.3 0.1 ;
  LAYER metal5 ;
        RECT -0.56 -0.1 0.16  0.1 ;
END VIA45_DC_LEFT

VIA VIA45_DC_TOP DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.16 0.1 0.56 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 0.3 0.1 0.5 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.16  0.5 ;
END VIA45_DC_TOP

VIA VIA45_DC_DOWN DEFAULT
  LAYER metal4 ;
        RECT -0.1 -0.56 0.1 0.16 ;
  LAYER via4 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 -0.5 0.1 -0.3 ;
  LAYER metal5 ;
        RECT -0.16 -0.5 0.16  0.1 ;
END VIA45_DC_DOWN

VIA VIA56_DC_RIGHT DEFAULT
  LAYER metal6 ;
        RECT -0.1 -0.16 0.5 0.16 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT 0.3 -0.1 0.5 0.1 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.56  0.1 ;
END VIA56_DC_RIGHT

VIA VIA56_DC_LEFT DEFAULT
  LAYER metal6 ;
        RECT -0.5 -0.16 0.1 0.16 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.5 -0.1 -0.3 0.1 ;
  LAYER metal5 ;
        RECT -0.56 -0.1 0.16  0.1 ;
END VIA56_DC_LEFT

VIA VIA56_DC_TOP DEFAULT
  LAYER metal6 ;
        RECT -0.1 -0.16 0.1 0.56 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 0.3 0.1 0.5 ;
  LAYER metal5 ;
        RECT -0.16 -0.1 0.16  0.5 ;
END VIA56_DC_TOP

VIA VIA56_DC_DOWN DEFAULT
  LAYER metal6 ;
        RECT -0.1 -0.56 0.1 0.16 ;
  LAYER via5 ;
        RECT -0.1 -0.1 0.1 0.1 ;
        RECT -0.1 -0.5 0.1 -0.3 ;
  LAYER metal5 ;
        RECT -0.16 -0.5 0.16  0.1 ;
END VIA56_DC_DOWN

VIA VIA67_DC_RIGHT DEFAULT
  LAYER metal6 ;
        RECT -0.2 -0.2 1.0 0.2 ;
  LAYER via6 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT 0.6 -0.2 1.0 0.2 ;
  LAYER metal7 ;
        RECT -0.2 -0.2 1.0  0.2 ;
END VIA67_DC_RIGHT

VIA VIA67_DC_LEFT DEFAULT
  LAYER metal6 ;
        RECT -1.0 -0.2 0.2 0.2 ;
  LAYER via6 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT -1.0 -0.2 -0.6 0.2 ;
  LAYER metal7 ;
        RECT -1.0 -0.2 0.2  0.2 ;
END VIA67_DC_LEFT

VIA VIA67_DC_TOP DEFAULT
  LAYER metal6 ;
        RECT -0.2 -0.2 0.2 1.0 ;
  LAYER via6 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT -0.2 0.6 0.2 1.0 ;
  LAYER metal7 ;
        RECT -0.2 -0.2 0.2  1.0 ;
END VIA67_DC_TOP

VIA VIA67_DC_DOWN DEFAULT
  LAYER metal6 ;
        RECT -0.2 -1.0 0.2 0.2 ;
  LAYER via6 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT -0.2 -1.0 0.2 -0.6 ;
  LAYER metal7 ;
        RECT -0.2 -1.0 0.2  0.2 ;
END VIA67_DC_DOWN

VIA VIA78_DC_RIGHT DEFAULT
  LAYER metal8 ;
        RECT -0.2 -0.2 1.0 0.2 ;
  LAYER via7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT 0.6 -0.2 1.0 0.2 ;
  LAYER metal7 ;
        RECT -0.2 -0.2 1.0  0.2 ;
END VIA78_DC_RIGHT

VIA VIA78_DC_LEFT DEFAULT
  LAYER metal8 ;
        RECT -1.0 -0.2 0.2 0.2 ;
  LAYER via7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT -1.0 -0.2 -0.6 0.2 ;
  LAYER metal7 ;
        RECT -1.0 -0.2 0.2  0.2 ;
END VIA78_DC_LEFT

VIA VIA78_DC_TOP DEFAULT
  LAYER metal8 ;
        RECT -0.2 -0.2 0.2 1.0 ;
  LAYER via7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT -0.2 0.6 0.2 1.0 ;
  LAYER metal7 ;
        RECT -0.2 -0.2 0.2  1.0 ;
END VIA78_DC_TOP

VIA VIA78_DC_DOWN DEFAULT
  LAYER metal8 ;
        RECT -0.2 -1.0 0.2 0.2 ;
  LAYER via7 ;
        RECT -0.2 -0.2 0.2 0.2 ;
        RECT -0.2 -1.0 0.2 -0.6 ;
  LAYER metal7 ;
        RECT -0.2 -1.0 0.2  0.2 ;
END VIA78_DC_DOWN

#------------------------------------------


#------------------------------------------
# define via rules for via usage
# while invoking SROUTE, ADD WIRE, or MOVE WIRE command
#------------------------------------------

# vias generated from signal via rules

VIA VIA12_HH_2cut_E DEFAULT 
    LAYER metal1 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
END VIA12_HH_2cut_E
VIA VIA12_HH_2cut_W DEFAULT 
    LAYER metal1 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal2 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
END VIA12_HH_2cut_W
VIA VIA12_HH_2cut_N DEFAULT 
    LAYER metal1 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    LAYER via ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
END VIA12_HH_2cut_N
VIA VIA12_HH_2cut_S DEFAULT 
    LAYER metal1 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    LAYER via ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal2 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
END VIA12_HH_2cut_S
VIA VIA12_HH_2cut_alt_E DEFAULT 
    LAYER metal1 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
END VIA12_HH_2cut_alt_E
VIA VIA12_HH_2cut_alt_W DEFAULT 
    LAYER metal1 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal2 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
END VIA12_HH_2cut_alt_W
VIA VIA12_HH_2cut_alt_N DEFAULT 
    LAYER metal1 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    LAYER via ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal2 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
END VIA12_HH_2cut_alt_N
VIA VIA12_HH_2cut_alt_S DEFAULT 
    LAYER metal1 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    LAYER via ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal2 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
END VIA12_HH_2cut_alt_S
VIA VIA23_HH_mar_N DEFAULT  TOPOFSTACKONLY
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.160000 0.220000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA23_HH_mar_N
VIA VIA23_HH_mar_S DEFAULT  TOPOFSTACKONLY
    LAYER metal2 ; 
	RECT -0.160000 -0.220000 0.160000 0.100000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA23_HH_mar_S
VIA VIA23_HH_2cut_E DEFAULT 
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_E
VIA VIA23_HH_2cut_W DEFAULT 
    LAYER metal2 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via2 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_W
VIA VIA23_HH_2cut_N DEFAULT 
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_N
VIA VIA23_HH_2cut_S DEFAULT 
    LAYER metal2 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_S
VIA VIA23_HH_2cut_alt_E DEFAULT 
    LAYER metal2 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_alt_E
VIA VIA23_HH_2cut_alt_W DEFAULT 
    LAYER metal2 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via2 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_alt_W
VIA VIA23_HH_2cut_alt_N DEFAULT 
    LAYER metal2 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal3 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_alt_N
VIA VIA23_HH_2cut_alt_S DEFAULT 
    LAYER metal2 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    LAYER via2 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal3 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    RESISTANCE 0.750000 ;
END VIA23_HH_2cut_alt_S
VIA VIA34_HH_mar_E DEFAULT  TOPOFSTACKONLY
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.360000 0.100000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA34_HH_mar_E
VIA VIA34_HH_mar_W DEFAULT  TOPOFSTACKONLY
    LAYER metal3 ; 
	RECT -0.360000 -0.100000 0.160000 0.100000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA34_HH_mar_W
VIA VIA34_HH_2cut_E DEFAULT 
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_E
VIA VIA34_HH_2cut_W DEFAULT 
    LAYER metal3 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via3 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_W
VIA VIA34_HH_2cut_N DEFAULT 
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_N
VIA VIA34_HH_2cut_S DEFAULT 
    LAYER metal3 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_S
VIA VIA34_HH_2cut_alt_E DEFAULT 
    LAYER metal3 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_alt_E
VIA VIA34_HH_2cut_alt_W DEFAULT 
    LAYER metal3 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via3 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_alt_W
VIA VIA34_HH_2cut_alt_N DEFAULT 
    LAYER metal3 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal4 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_alt_N
VIA VIA34_HH_2cut_alt_S DEFAULT 
    LAYER metal3 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    LAYER via3 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal4 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    RESISTANCE 0.750000 ;
END VIA34_HH_2cut_alt_S
VIA VIA45_HH_mar_N DEFAULT  TOPOFSTACKONLY
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.160000 0.220000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA45_HH_mar_N
VIA VIA45_HH_mar_S DEFAULT  TOPOFSTACKONLY
    LAYER metal4 ; 
	RECT -0.160000 -0.220000 0.160000 0.100000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA45_HH_mar_S
VIA VIA45_HH_2cut_E DEFAULT 
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_E
VIA VIA45_HH_2cut_W DEFAULT 
    LAYER metal4 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via4 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_W
VIA VIA45_HH_2cut_N DEFAULT 
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_N
VIA VIA45_HH_2cut_S DEFAULT 
    LAYER metal4 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_S
VIA VIA45_HH_2cut_alt_E DEFAULT 
    LAYER metal4 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_alt_E
VIA VIA45_HH_2cut_alt_W DEFAULT 
    LAYER metal4 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via4 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_alt_W
VIA VIA45_HH_2cut_alt_N DEFAULT 
    LAYER metal4 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal5 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_alt_N
VIA VIA45_HH_2cut_alt_S DEFAULT 
    LAYER metal4 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    LAYER via4 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal5 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    RESISTANCE 0.750000 ;
END VIA45_HH_2cut_alt_S
VIA VIA56_HH_mar_E DEFAULT  TOPOFSTACKONLY
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.360000 0.100000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA56_HH_mar_E
VIA VIA56_HH_mar_W DEFAULT  TOPOFSTACKONLY
    LAYER metal5 ; 
	RECT -0.360000 -0.100000 0.160000 0.100000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.160000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 1.500000 ;
END VIA56_HH_mar_W
VIA VIA56_HH_2cut_E DEFAULT 
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_E
VIA VIA56_HH_2cut_W DEFAULT 
    LAYER metal5 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via5 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_W
VIA VIA56_HH_2cut_N DEFAULT 
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal6 ; 
	RECT -0.160000 -0.100000 0.160000 0.500000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_N
VIA VIA56_HH_2cut_S DEFAULT 
    LAYER metal5 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.160000 -0.500000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_S
VIA VIA56_HH_2cut_alt_E DEFAULT 
    LAYER metal5 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT 0.300000 -0.100000 0.500000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.160000 -0.100000 0.560000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_alt_E
VIA VIA56_HH_2cut_alt_W DEFAULT 
    LAYER metal5 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    LAYER via5 ; 
	RECT -0.500000 -0.100000 -0.300000 0.100000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.560000 -0.100000 0.160000 0.100000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_alt_W
VIA VIA56_HH_2cut_alt_N DEFAULT 
    LAYER metal5 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
	RECT -0.100000 0.300000 0.100000 0.500000 ;
    LAYER metal6 ; 
	RECT -0.100000 -0.160000 0.100000 0.560000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_alt_N
VIA VIA56_HH_2cut_alt_S DEFAULT 
    LAYER metal5 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    LAYER via5 ; 
	RECT -0.100000 -0.500000 0.100000 -0.300000 ;
	RECT -0.100000 -0.100000 0.100000 0.100000 ;
    LAYER metal6 ; 
	RECT -0.100000 -0.560000 0.100000 0.160000 ;
    RESISTANCE 0.750000 ;
END VIA56_HH_2cut_alt_S

# end auto generated vias

VIARULE VIAM1M2A
   LAYER metal1 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.160 to 0.160 ;
   LAYER metal2 ;
      DIRECTION VERTICAL ;
      WIDTH 0.200 to 0.200 ;
   VIA VIA12_HH ;
   VIA VIA12_VH ;
   VIA VIA12_HV ;
   VIA VIA12_VV ;
END VIAM1M2A

VIARULE VIAM2M3
   LAYER metal2 ;
      DIRECTION VERTICAL ;
      WIDTH 0.200 to 0.200 ;
   LAYER metal3 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.200 to 0.200 ;
   VIA VIA23_HH ;
   VIA VIA23_VH ;
   VIA VIA23_HV ;
   VIA VIA23_VV ;
END VIAM2M3

VIARULE VIAM3M4
   LAYER metal3 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.200 to 0.200 ;
   LAYER metal4 ;
      DIRECTION VERTICAL ;
      WIDTH 0.200 to 0.200 ;
   VIA VIA34_HH ;
   VIA VIA34_VH ;
   VIA VIA34_HV ;
   VIA VIA34_VV ;
END VIAM3M4

VIARULE VIAM4M5
   LAYER metal4 ;
      DIRECTION VERTICAL ;
      WIDTH 0.200 to 0.200 ;
   LAYER metal5 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.200 to 0.200 ;
   VIA VIA45_HH ;
   VIA VIA45_VH ;
   VIA VIA45_HV ;
   VIA VIA45_VV ;
END VIAM4M5

VIARULE VIAM5M6
   LAYER metal5 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.200 to 0.200 ;
   LAYER metal6 ;
      DIRECTION VERTICAL ;
      WIDTH 0.200 to 0.200 ;
   VIA VIA56_HH ;
   VIA VIA56_VH ;
   VIA VIA56_HV ;
   VIA VIA56_VV ;
END VIAM5M6

VIARULE VIAM6M7
   LAYER metal6 ;
      DIRECTION VERTICAL ;
      WIDTH 0.200 to 0.200 ;
   LAYER metal7 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.400 to 0.400 ;
   VIA VIA67_Def ;
END VIAM6M7
 
VIARULE VIAM7M8
   LAYER metal7 ;
      DIRECTION HORIZONTAL ;
      WIDTH 0.400 to 0.400 ;
   LAYER metal8 ;
      DIRECTION VERTICAL ;
      WIDTH 0.400 to 0.400 ;
   VIA VIA78_Def ;
END VIAM7M8

#------------------------------------------
# turn via rules fill in the corner area at the intersection
# between two speial wires at the same layer, where each wire
# must be extended by half the width of the other wire.
#------------------------------------------

#viarule turn1 generate
#   layer metal1 ;
#   direction horizontal ;
#   layer metal1 ;
#   direction vertical ;
#end turn1

#viarule turn2 generate
#   layer metal2 ;
#   direction horizontal ;
#   layer metal2 ;
#   direction vertical ;
#end turn2

#viarule turn3 generate
#   layer metal3 ;
#   direction horizontal ;
#   layer metal3 ;
#   direction vertical ;
#end turn3

#viarule turn4 generate
#   layer metal4 ;
#   direction horizontal ;
#   layer metal4 ;
#   direction vertical ;
#end turn4

#viarule turn5 generate
#   layer metal5 ;
#   direction horizontal ;
#   layer metal5 ;
#   direction vertical ;
#end turn5

#viarule turn6 generate
#   layer metal6 ;
#   direction horizontal ;
#   layer metal6 ;
#   direction vertical ;
#end turn6

#viarule turn7 generate
#   layer metal7 ;
#   direction horizontal ;
#   layer metal7 ;
#   direction vertical ;
#end turn7

#viarule turn8 generate
#   layer metal8 ;
#   direction horizontal ;
#   layer metal8 ;
#   direction vertical ;
#end turn8

#------------------------------------------
# define the a formula of via array generation 1
#------------------------------------------
viarule genm1m2a generate
   layer metal1 ;
      direction horizontal ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal2 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm1m2a

viarule genm1m2b generate
   layer metal1 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal2 ;
      direction vertical ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm1m2b


viarule genm2m3a generate
   layer metal2 ;
      direction vertical ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal3 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via2 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm2m3a

viarule genm2m3b generate
   layer metal2 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal3 ;
      direction horizontal ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via2 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm2m3b

viarule genm3m4a generate
   layer metal3 ;
      direction horizontal ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal4 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via3 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm3m4a

viarule genm3m4b generate
   layer metal3 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal4 ;
      direction vertical ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via3 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm3m4b


viarule genm4m5a generate
   layer metal4 ;
      direction vertical ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal5 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via4 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm4m5a

viarule genm4m5b generate
   layer metal4 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal5 ;
      direction horizontal ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via4 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm4m5b

viarule genm5m6a generate
   layer metal5 ;
      direction horizontal ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal6 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via5 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm5m6a

viarule genm5m6b generate
   layer metal5 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal6 ;
      direction vertical ;
      width 0.01 to 1.11 ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via5 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.400 by 0.400 ;
end genm5m6b

viarule genm6m7a generate
   layer metal6 ;
      direction vertical ;
      width 0.01 to 1.99 ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer metal7 ;
      direction horizontal ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer via6 ;
      rect -0.200 -0.200 0.200 0.200 ;
      spacing 0.800 by 0.800 ;
end genm6m7a
 
viarule genm6m7b generate
   layer metal6 ;
      direction vertical ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer metal7 ;
      direction horizontal ;
      width 0.01 to 1.99 ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer via6 ;
      rect -0.200 -0.200 0.200 0.200 ;
      spacing 0.800 by 0.800 ;
end genm6m7b

viarule genm7m8a generate
   layer metal7 ;
      direction horizontal ;
      width 0.01 to 1.99 ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer metal8 ;
      direction vertical ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer via7 ;
      rect -0.200 -0.200 0.200 0.200 ;
      spacing 0.800 by 0.800 ;
end genm7m8a

viarule genm7m8b generate
   layer metal7 ;
      direction horizontal ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer metal8 ;
      direction vertical ;
      width 0.01 to 1.99 ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer via7 ;
      rect -0.200 -0.200 0.200 0.200 ;
      spacing 0.800 by 0.800 ;
end genm7m8b


#------------------------------------------
# define the a formula of via array generation 2 for array >= 3x3
#------------------------------------------
viarule genm1m2_w generate
   layer metal1 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal2 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.480 by 0.480 ;
end genm1m2_w

viarule genm2m3_w generate
   layer metal2 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal3 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via2 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.480 by 0.480 ;
end genm2m3_w

viarule genm3m4_w generate
   layer metal3 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal4 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via3 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.480 by 0.480 ;
end genm3m4_w

viarule genm4m5_w generate
   layer metal4 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal5 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via4 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.480 by 0.480 ;
end genm4m5_w

viarule genm5m6_w generate
   layer metal5 ;
      direction horizontal ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer metal6 ;
      direction vertical ;
      overhang .060 ;
      metaloverhang 0.0 ;
   layer via5 ;
      rect -0.100 -0.100 0.100 0.100 ;
      spacing 0.480 by 0.480 ;
end genm5m6_w

viarule genm6m7_w generate
   layer metal6 ;
      direction vertical ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer metal7 ;
      direction horizontal ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer via6 ;
      rect -0.200 -0.200 0.200 0.200 ;
      spacing 0.900 by 0.900 ;
end genm6m7_w
 
viarule genm7m8_w generate
   layer metal7 ;
      direction horizontal ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer metal8 ;
      direction vertical ;
      overhang .000 ;
      metaloverhang 0.0 ;
   layer via7 ;
      rect -0.200 -0.200 0.200 0.200 ;
      spacing 0.900 by 0.900 ;
end genm7m8_w

#------------------------------------------
# define the samenet spacing table gives the samenet
# spacing rule
#------------------------------------------
#SPACING
#   SAMENET contact via 0 stack ;
#   SAMENET metal1 metal1 0.16 stack ;
#   SAMENET via via 0.20 ;
#   SAMENET metal2 metal2 0.20 stack ;
#   SAMENET via via2 0 stack ;
#   SAMENET via2 via2 0.20 ;
#   SAMENET metal3 metal3 0.20 stack ;
#   SAMENET via2 via3 0 stack ;
#   SAMENET via3 via3 0.20 ;
#   SAMENET metal4 metal4 0.20 stack ;
#   SAMENET via3 via4 0 stack ;
#   SAMENET via4 via4 0.20 ;
#   SAMENET metal5 metal5 0.20 stack ;
#   SAMENET via4 via5 0 stack ;
#   SAMENET via5 via5 0.20 ;
#   SAMENET metal6 metal6 0.20 stack ;
#   SAMENET via5 via6 0 stack ;
#   SAMENET via6 via6 0.40 ;
#   SAMENET metal7 metal7 0.40 stack ;
#   SAMENET via6 via7 0 stack ;
#   SAMENET via7 via7 0.40 ;
#   SAMENET metal8 metal8 0.40 ;
#END SPACING

#------------------------------------------
# site definition for P&R
#------------------------------------------
SITE core
    SYMMETRY y ;
    CLASS CORE  ;
    SIZE 0.400 BY 3.200 ;
END core

SITE core_3200
    SYMMETRY y ;
    CLASS CORE  ;
    SIZE 0.400 BY 3.200 ;
END core_3200

SITE core_2800
    SYMMETRY y ;
    CLASS CORE  ;
    SIZE 0.400 BY 2.800 ;
END core_2800

SITE corega_3200
    SYMMETRY y ;
    CLASS CORE  ;
    SIZE 2.00 BY 3.20 ;
END corega_3200

SITE iocore_a
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 218.400 ;
END iocore_a

SITE iocore_b
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 152.000 ;
END iocore_b

SITE iocore_as
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 242.800 ;
END iocore_as

SITE iocore_bs
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 169.200 ;
END iocore_bs

SITE iocore_k
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 268.000 ;
END iocore_k

SITE iocore_n
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 282.800 ;
END iocore_n

SITE iocore_o
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 206.00 ;
END iocore_o

SITE corner_a
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 218.400 BY 218.400 ;
END corner_a

SITE corner_b
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 152.000 BY 152.000 ;
END corner_b

SITE corner_ab
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 218.400 BY 152.000 ;
END corner_ab

SITE iocore_c
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 172.00 ;
END iocore_c

SITE iocore_d
    SYMMETRY y ;
    CLASS PAD  ;
    SIZE 0.400 BY 104.00 ;
END iocore_d


END LIBRARY
