##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Wed Dec 15 19:38:08 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERbg
  CLASS BLOCK ;
  SIZE 120.000000 BY 40.000000 ;
  FOREIGN BATCHARGERbg 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 20.120000 39.360000 20.280000 40.000000 ;
    END
  END vin
  PIN ibias1ua
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 2.120000 0.640000 2.280000 ;
    END
  END ibias1ua
  PIN ibias1ub
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 0.120000 0.640000 0.280000 ;
    END
  END ibias1ub
  PIN vrefa
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 4.120000 0.640000 4.280000 ;
    END
  END vrefa
  PIN vrefb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 6.120000 0.640000 6.280000 ;
    END
  END vrefb
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.120000 39.360000 10.280000 40.000000 ;
    END
  END en
  PIN endvdd
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.120000 39.360000 12.280000 40.000000 ;
    END
  END endvdd
  PIN clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.120000 39.360000 4.280000 40.000000 ;
    END
  END clk
  PIN rstz
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.120000 39.360000 18.280000 40.000000 ;
    END
  END rstz
  PIN avdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 110.500000 0.000000 111.500000 0.640000 ;
    END
  END avdd
  PIN dvdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 100.500000 0.000000 101.500000 0.640000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 100.500000 39.360000 101.500000 40.000000 ;
    END
  END dgnd
  PIN agnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 110.500000 39.360000 111.500000 40.000000 ;
    END
  END agnd
  OBS
    LAYER metal1 ;
      RECT 111.660000 39.200000 120.000000 40.000000 ;
      RECT 101.660000 39.200000 110.340000 40.000000 ;
      RECT 20.440000 39.200000 100.340000 40.000000 ;
      RECT 18.440000 39.200000 19.960000 40.000000 ;
      RECT 12.440000 39.200000 17.960000 40.000000 ;
      RECT 10.440000 39.200000 11.960000 40.000000 ;
      RECT 4.440000 39.200000 9.960000 40.000000 ;
      RECT 0.000000 39.200000 3.960000 40.000000 ;
      RECT 0.000000 6.440000 120.000000 39.200000 ;
      RECT 0.830000 5.960000 120.000000 6.440000 ;
      RECT 0.000000 4.440000 120.000000 5.960000 ;
      RECT 0.830000 3.960000 120.000000 4.440000 ;
      RECT 0.000000 2.440000 120.000000 3.960000 ;
      RECT 0.830000 1.960000 120.000000 2.440000 ;
      RECT 0.000000 0.800000 120.000000 1.960000 ;
      RECT 0.000000 0.440000 100.340000 0.800000 ;
      RECT 111.660000 0.000000 120.000000 0.800000 ;
      RECT 101.660000 0.000000 110.340000 0.800000 ;
      RECT 0.830000 0.000000 100.340000 0.440000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
    LAYER metal3 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 120.000000 40.000000 ;
  END
END BATCHARGERbg

END LIBRARY
