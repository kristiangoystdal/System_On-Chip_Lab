VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO GNDACUTHA
    CLASS PAD ;
    FOREIGN GNDACUTHA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.200 BY 218.400 ;
    SYMMETRY x y r90 ;
    SITE iocore_a ;
    PIN GNDANA
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal7 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal6 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal5 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal4 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal3 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal2 ;
        RECT  13.860 213.450 23.600 218.000 ;
        LAYER metal1 ;
        RECT  13.860 213.450 23.600 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal7 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal6 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal5 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal4 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal3 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal2 ;
        RECT  1.600 213.450 11.340 218.000 ;
        LAYER metal1 ;
        RECT  1.600 213.450 11.340 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal7 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal6 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal5 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal4 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal3 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal2 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal1 ;
        RECT  1.600 0.000 23.600 3.480 ;
        END
    END GNDANA
    OBS
        LAYER metal1 ;
        POLYGON  25.200 217.800 23.860 217.800 23.860 213.190 13.600 213.190
                 13.600 217.800 11.600 217.800 11.600 213.190 1.340 213.190 1.340 217.800
                 0.000 217.800 0.000 0.000 1.340 0.000 1.340 3.740 23.860 3.740
                 23.860 0.000 25.200 0.000 ;
        LAYER via ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal2 ;
        POLYGON  25.200 217.800 23.880 217.800 23.880 213.170 13.580 213.170
                 13.580 217.800 11.620 217.800 11.620 213.170 1.320 213.170 1.320 217.800
                 0.000 217.800 0.000 0.000 1.320 0.000 1.320 3.760 23.880 3.760
                 23.880 0.000 25.200 0.000 ;
        LAYER via2 ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal3 ;
        POLYGON  25.200 217.800 23.880 217.800 23.880 213.170 13.580 213.170
                 13.580 217.800 11.620 217.800 11.620 213.170 1.320 213.170 1.320 217.800
                 0.000 217.800 0.000 0.000 1.320 0.000 1.320 3.760 23.880 3.760
                 23.880 0.000 25.200 0.000 ;
        LAYER via3 ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal4 ;
        POLYGON  25.200 217.800 23.880 217.800 23.880 213.170 13.580 213.170
                 13.580 217.800 11.620 217.800 11.620 213.170 1.320 213.170 1.320 217.800
                 0.000 217.800 0.000 0.000 1.320 0.000 1.320 3.760 23.880 3.760
                 23.880 0.000 25.200 0.000 ;
        LAYER via4 ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal5 ;
        POLYGON  25.200 217.800 24.100 217.800 24.100 212.950 13.360 212.950
                 13.360 217.800 11.840 217.800 11.840 212.950 1.100 212.950 1.100 217.800
                 0.000 217.800 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
        LAYER via5 ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal6 ;
        POLYGON  25.200 217.800 24.100 217.800 24.100 212.950 13.360 212.950
                 13.360 217.800 11.840 217.800 11.840 212.950 1.100 212.950 1.100 217.800
                 0.000 217.800 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
        LAYER via6 ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal7 ;
        POLYGON  25.200 217.800 24.100 217.800 24.100 212.950 13.360 212.950
                 13.360 217.800 11.840 217.800 11.840 212.950 1.100 212.950 1.100 217.800
                 0.000 217.800 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
        LAYER via7 ;
        RECT  13.860 213.450 23.600 218.000 ;
        RECT  1.600 213.450 11.340 218.000 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal8 ;
        POLYGON  25.200 217.800 24.100 217.800 24.100 212.950 13.360 212.950
                 13.360 217.800 11.840 217.800 11.840 212.950 1.100 212.950 1.100 217.800
                 0.000 217.800 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
    END
END GNDACUTHA

MACRO GNDACUTHB
    CLASS PAD ;
    FOREIGN GNDACUTHB 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.200 BY 152.000 ;
    SYMMETRY x y r90 ;
    SITE iocore_b ;
    PIN GNDANA
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal7 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal6 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal5 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal4 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal3 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal2 ;
        RECT  13.860 147.050 23.600 151.600 ;
        LAYER metal1 ;
        RECT  13.860 147.050 23.600 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal7 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal6 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal5 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal4 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal3 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal2 ;
        RECT  1.600 147.050 11.340 151.600 ;
        LAYER metal1 ;
        RECT  1.600 147.050 11.340 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal7 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal6 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal5 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal4 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal3 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal2 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal1 ;
        RECT  1.600 0.000 23.600 3.480 ;
        END
    END GNDANA
    OBS
        LAYER metal1 ;
        POLYGON  25.200 151.400 23.860 151.400 23.860 146.790 13.600 146.790
                 13.600 151.400 11.600 151.400 11.600 146.790 1.340 146.790 1.340 151.400
                 0.000 151.400 0.000 0.000 1.340 0.000 1.340 3.740 23.860 3.740
                 23.860 0.000 25.200 0.000 ;
        LAYER via ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal2 ;
        POLYGON  25.200 151.400 23.880 151.400 23.880 146.770 13.580 146.770
                 13.580 151.400 11.620 151.400 11.620 146.770 1.320 146.770 1.320 151.400
                 0.000 151.400 0.000 0.000 1.320 0.000 1.320 3.760 23.880 3.760
                 23.880 0.000 25.200 0.000 ;
        LAYER via2 ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal3 ;
        POLYGON  25.200 151.400 23.880 151.400 23.880 146.770 13.580 146.770
                 13.580 151.400 11.620 151.400 11.620 146.770 1.320 146.770 1.320 151.400
                 0.000 151.400 0.000 0.000 1.320 0.000 1.320 3.760 23.880 3.760
                 23.880 0.000 25.200 0.000 ;
        LAYER via3 ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal4 ;
        POLYGON  25.200 151.400 23.880 151.400 23.880 146.770 13.580 146.770
                 13.580 151.400 11.620 151.400 11.620 146.770 1.320 146.770 1.320 151.400
                 0.000 151.400 0.000 0.000 1.320 0.000 1.320 3.760 23.880 3.760
                 23.880 0.000 25.200 0.000 ;
        LAYER via4 ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal5 ;
        POLYGON  25.200 151.400 24.100 151.400 24.100 146.550 13.360 146.550
                 13.360 151.400 11.840 151.400 11.840 146.550 1.100 146.550 1.100 151.400
                 0.000 151.400 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
        LAYER via5 ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal6 ;
        POLYGON  25.200 151.400 24.100 151.400 24.100 146.550 13.360 146.550
                 13.360 151.400 11.840 151.400 11.840 146.550 1.100 146.550 1.100 151.400
                 0.000 151.400 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
        LAYER via6 ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal7 ;
        POLYGON  25.200 151.400 24.100 151.400 24.100 146.550 13.360 146.550
                 13.360 151.400 11.840 151.400 11.840 146.550 1.100 146.550 1.100 151.400
                 0.000 151.400 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
        LAYER via7 ;
        RECT  13.860 147.050 23.600 151.600 ;
        RECT  1.600 147.050 11.340 151.600 ;
        RECT  1.600 0.000 23.600 3.480 ;
        LAYER metal8 ;
        POLYGON  25.200 151.400 24.100 151.400 24.100 146.550 13.360 146.550
                 13.360 151.400 11.840 151.400 11.840 146.550 1.100 146.550 1.100 151.400
                 0.000 151.400 0.000 0.000 1.100 0.000 1.100 3.980 24.100 3.980
                 24.100 0.000 25.200 0.000 ;
    END
END GNDACUTHB

MACRO LCUT12HA
    CLASS PAD ;
    FOREIGN LCUT12HA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 48.000 BY 218.400 ;
    SYMMETRY x y r90 ;
    SITE iocore_a ;
    PIN VCC12VESD
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal7 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal6 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal5 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal4 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal3 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal2 ;
        RECT  9.720 213.450 25.920 218.000 ;
        LAYER metal1 ;
        RECT  9.720 213.450 25.920 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal7 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal6 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal5 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal4 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal3 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal2 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal1 ;
        RECT  29.280 213.450 45.480 218.000 ;
        END
    END VCC12VESD
    OBS
        LAYER metal1 ;
        POLYGON  48.000 218.000 45.740 218.000 45.740 213.190 29.020 213.190
                 29.020 218.000 26.180 218.000 26.180 213.190 9.460 213.190 9.460 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal2 ;
        POLYGON  48.000 218.000 45.760 218.000 45.760 213.170 29.000 213.170
                 29.000 218.000 26.200 218.000 26.200 213.170 9.440 213.170 9.440 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via2 ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal3 ;
        POLYGON  48.000 218.000 45.760 218.000 45.760 213.170 29.000 213.170
                 29.000 218.000 26.200 218.000 26.200 213.170 9.440 213.170 9.440 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via3 ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal4 ;
        POLYGON  48.000 218.000 45.760 218.000 45.760 213.170 29.000 213.170
                 29.000 218.000 26.200 218.000 26.200 213.170 9.440 213.170 9.440 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via4 ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal5 ;
        POLYGON  48.000 218.000 45.980 218.000 45.980 212.950 28.780 212.950
                 28.780 218.000 26.420 218.000 26.420 212.950 9.220 212.950 9.220 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via5 ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal6 ;
        POLYGON  48.000 218.000 45.980 218.000 45.980 212.950 28.780 212.950
                 28.780 218.000 26.420 218.000 26.420 212.950 9.220 212.950 9.220 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via6 ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal7 ;
        POLYGON  48.000 218.000 45.980 218.000 45.980 212.950 28.780 212.950
                 28.780 218.000 26.420 218.000 26.420 212.950 9.220 212.950 9.220 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
        LAYER via7 ;
        RECT  9.720 213.450 25.920 218.000 ;
        RECT  29.280 213.450 45.480 218.000 ;
        LAYER metal8 ;
        POLYGON  48.000 218.000 45.980 218.000 45.980 212.950 28.780 212.950
                 28.780 218.000 26.420 218.000 26.420 212.950 9.220 212.950 9.220 218.000
                 0.000 218.000 0.000 0.000 48.000 0.000 ;
    END
END LCUT12HA

MACRO LCUT12HB
    CLASS PAD ;
    FOREIGN LCUT12HB 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 69.200 BY 152.000 ;
    SYMMETRY x y r90 ;
    SITE iocore_b ;
    PIN VCC12VESD
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal7 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal6 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal5 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal4 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal3 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal2 ;
        RECT  39.880 147.050 64.360 151.600 ;
        LAYER metal1 ;
        RECT  39.880 147.050 64.360 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal7 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal6 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal5 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal4 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal3 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal2 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal1 ;
        RECT  12.040 147.050 36.520 151.600 ;
        END
    END VCC12VESD
    OBS
        LAYER metal1 ;
        POLYGON  69.200 151.600 64.620 151.600 64.620 146.790 39.620 146.790
                 39.620 151.600 36.780 151.600 36.780 146.790 11.780 146.790
                 11.780 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal2 ;
        POLYGON  69.200 151.600 64.640 151.600 64.640 146.770 39.600 146.770
                 39.600 151.600 36.800 151.600 36.800 146.770 11.760 146.770
                 11.760 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via2 ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal3 ;
        POLYGON  69.200 151.600 64.640 151.600 64.640 146.770 39.600 146.770
                 39.600 151.600 36.800 151.600 36.800 146.770 11.760 146.770
                 11.760 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via3 ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal4 ;
        POLYGON  69.200 151.600 64.640 151.600 64.640 146.770 39.600 146.770
                 39.600 151.600 36.800 151.600 36.800 146.770 11.760 146.770
                 11.760 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via4 ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal5 ;
        POLYGON  69.200 151.600 64.860 151.600 64.860 146.550 39.380 146.550
                 39.380 151.600 37.020 151.600 37.020 146.550 11.540 146.550
                 11.540 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via5 ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal6 ;
        POLYGON  69.200 151.600 64.860 151.600 64.860 146.550 39.380 146.550
                 39.380 151.600 37.020 151.600 37.020 146.550 11.540 146.550
                 11.540 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via6 ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal7 ;
        POLYGON  69.200 151.600 64.860 151.600 64.860 146.550 39.380 146.550
                 39.380 151.600 37.020 151.600 37.020 146.550 11.540 146.550
                 11.540 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
        LAYER via7 ;
        RECT  39.880 147.050 64.360 151.600 ;
        RECT  12.040 147.050 36.520 151.600 ;
        LAYER metal8 ;
        POLYGON  69.200 151.600 64.860 151.600 64.860 146.550 39.380 146.550
                 39.380 151.600 37.020 151.600 37.020 146.550 11.540 146.550
                 11.540 151.600 0.000 151.600 0.000 0.000 69.200 0.000 ;
    END
END LCUT12HB

MACRO RCUT12HA
    CLASS PAD ;
    FOREIGN RCUT12HA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 57.200 BY 218.400 ;
    SYMMETRY x y r90 ;
    SITE iocore_a ;
    PIN GNDVESD
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal7 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal6 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal5 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal4 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal3 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal2 ;
        RECT  18.900 213.450 35.120 218.000 ;
        LAYER metal1 ;
        RECT  18.900 213.450 35.120 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal7 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal6 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal5 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal4 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal3 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal2 ;
        RECT  38.480 213.450 54.730 218.000 ;
        LAYER metal1 ;
        RECT  38.480 213.450 54.730 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal7 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal6 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal5 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal4 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal3 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal2 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal1 ;
        RECT  2.340 213.450 15.540 218.000 ;
        END
    END GNDVESD
    OBS
        LAYER metal1 ;
        POLYGON  57.200 218.000 54.990 218.000 54.990 213.190 38.220 213.190
                 38.220 218.000 35.380 218.000 35.380 213.190 18.640 213.190
                 18.640 218.000 15.800 218.000 15.800 213.190 2.080 213.190 2.080 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal2 ;
        POLYGON  57.200 218.000 55.010 218.000 55.010 213.170 38.200 213.170
                 38.200 218.000 35.400 218.000 35.400 213.170 18.620 213.170
                 18.620 218.000 15.820 218.000 15.820 213.170 2.060 213.170 2.060 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via2 ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal3 ;
        POLYGON  57.200 218.000 55.010 218.000 55.010 213.170 38.200 213.170
                 38.200 218.000 35.400 218.000 35.400 213.170 18.620 213.170
                 18.620 218.000 15.820 218.000 15.820 213.170 2.060 213.170 2.060 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via3 ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal4 ;
        POLYGON  57.200 218.000 55.010 218.000 55.010 213.170 38.200 213.170
                 38.200 218.000 35.400 218.000 35.400 213.170 18.620 213.170
                 18.620 218.000 15.820 218.000 15.820 213.170 2.060 213.170 2.060 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via4 ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal5 ;
        POLYGON  57.200 218.000 55.230 218.000 55.230 212.950 37.980 212.950
                 37.980 218.000 35.620 218.000 35.620 212.950 18.400 212.950
                 18.400 218.000 16.040 218.000 16.040 212.950 1.840 212.950 1.840 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via5 ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal6 ;
        POLYGON  57.200 218.000 55.230 218.000 55.230 212.950 37.980 212.950
                 37.980 218.000 35.620 218.000 35.620 212.950 18.400 212.950
                 18.400 218.000 16.040 218.000 16.040 212.950 1.840 212.950 1.840 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via6 ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal7 ;
        POLYGON  57.200 218.000 55.230 218.000 55.230 212.950 37.980 212.950
                 37.980 218.000 35.620 218.000 35.620 212.950 18.400 212.950
                 18.400 218.000 16.040 218.000 16.040 212.950 1.840 212.950 1.840 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
        LAYER via7 ;
        RECT  18.900 213.450 35.120 218.000 ;
        RECT  38.480 213.450 54.730 218.000 ;
        RECT  2.340 213.450 15.540 218.000 ;
        LAYER metal8 ;
        POLYGON  57.200 218.000 55.230 218.000 55.230 212.950 37.980 212.950
                 37.980 218.000 35.620 218.000 35.620 212.950 18.400 212.950
                 18.400 218.000 16.040 218.000 16.040 212.950 1.840 212.950 1.840 218.000
                 0.000 218.000 0.000 0.000 57.200 0.000 ;
    END
END RCUT12HA

MACRO RCUT12HB
    CLASS PAD ;
    FOREIGN RCUT12HB 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 82.400 BY 152.000 ;
    SYMMETRY x y r90 ;
    SITE iocore_b ;
    PIN GNDVESD
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal7 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal6 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal5 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal4 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal3 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal2 ;
        RECT  53.080 147.050 77.560 151.600 ;
        LAYER metal1 ;
        RECT  53.080 147.050 77.560 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal7 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal6 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal5 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal4 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal3 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal2 ;
        RECT  25.240 147.050 49.720 151.600 ;
        LAYER metal1 ;
        RECT  25.240 147.050 49.720 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal7 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal6 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal5 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal4 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal3 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal2 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal1 ;
        RECT  2.060 147.050 21.880 151.600 ;
        END
    END GNDVESD
    OBS
        LAYER metal1 ;
        POLYGON  82.400 151.600 77.820 151.600 77.820 146.790 52.820 146.790
                 52.820 151.600 49.980 151.600 49.980 146.790 24.980 146.790
                 24.980 151.600 22.140 151.600 22.140 146.790 1.800 146.790 1.800 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal2 ;
        POLYGON  82.400 151.600 77.840 151.600 77.840 146.770 52.800 146.770
                 52.800 151.600 50.000 151.600 50.000 146.770 24.960 146.770
                 24.960 151.600 22.160 151.600 22.160 146.770 1.780 146.770 1.780 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via2 ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal3 ;
        POLYGON  82.400 151.600 77.840 151.600 77.840 146.770 52.800 146.770
                 52.800 151.600 50.000 151.600 50.000 146.770 24.960 146.770
                 24.960 151.600 22.160 151.600 22.160 146.770 1.780 146.770 1.780 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via3 ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal4 ;
        POLYGON  82.400 151.600 77.840 151.600 77.840 146.770 52.800 146.770
                 52.800 151.600 50.000 151.600 50.000 146.770 24.960 146.770
                 24.960 151.600 22.160 151.600 22.160 146.770 1.780 146.770 1.780 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via4 ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal5 ;
        POLYGON  82.400 151.600 78.060 151.600 78.060 146.550 52.580 146.550
                 52.580 151.600 50.220 151.600 50.220 146.550 24.740 146.550
                 24.740 151.600 22.380 151.600 22.380 146.550 1.560 146.550 1.560 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via5 ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal6 ;
        POLYGON  82.400 151.600 78.060 151.600 78.060 146.550 52.580 146.550
                 52.580 151.600 50.220 151.600 50.220 146.550 24.740 146.550
                 24.740 151.600 22.380 151.600 22.380 146.550 1.560 146.550 1.560 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via6 ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal7 ;
        POLYGON  82.400 151.600 78.060 151.600 78.060 146.550 52.580 146.550
                 52.580 151.600 50.220 151.600 50.220 146.550 24.740 146.550
                 24.740 151.600 22.380 151.600 22.380 146.550 1.560 146.550 1.560 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
        LAYER via7 ;
        RECT  53.080 147.050 77.560 151.600 ;
        RECT  25.240 147.050 49.720 151.600 ;
        RECT  2.060 147.050 21.880 151.600 ;
        LAYER metal8 ;
        POLYGON  82.400 151.600 78.060 151.600 78.060 146.550 52.580 146.550
                 52.580 151.600 50.220 151.600 50.220 146.550 24.740 146.550
                 24.740 151.600 22.380 151.600 22.380 146.550 1.560 146.550 1.560 151.600
                 0.000 151.600 0.000 0.000 82.400 0.000 ;
    END
END RCUT12HB

MACRO ULSCI0CUTHA
    CLASS PAD ;
    FOREIGN ULSCI0CUTHA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.800 BY 218.400 ;
    SYMMETRY x y r90 ;
    SITE iocore_a ;
    PIN O
        DIRECTION INOUT ;
        PORT
        LAYER metal8 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal7 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal6 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal5 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal4 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal3 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal2 ;
        RECT  2.520 0.000 32.280 2.680 ;
        LAYER metal1 ;
        RECT  2.520 0.000 32.280 2.680 ;
        END
        PORT
        LAYER metal8 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal7 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal6 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal5 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal4 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal3 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal2 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal1 ;
        RECT  4.960 213.450 29.840 218.000 ;
        END
    END O
    PIN GNDANA
        DIRECTION INPUT ;
    END GNDANA
    PIN VCC12ANA
        DIRECTION INPUT ;
    END VCC12ANA
    OBS
        LAYER metal1 ;
        POLYGON  34.800 218.000 30.100 218.000 30.100 213.190 4.700 213.190 4.700 218.000
                 0.000 218.000 0.000 0.000 2.260 0.000 2.260 2.940 32.540 2.940
                 32.540 0.000 34.800 0.000 ;
        LAYER via ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal2 ;
        POLYGON  34.800 218.000 30.120 218.000 30.120 213.170 4.680 213.170 4.680 218.000
                 0.000 218.000 0.000 0.000 2.240 0.000 2.240 2.960 32.560 2.960
                 32.560 0.000 34.800 0.000 ;
        LAYER via2 ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal3 ;
        POLYGON  34.800 218.000 30.120 218.000 30.120 213.170 4.680 213.170 4.680 218.000
                 0.000 218.000 0.000 0.000 2.240 0.000 2.240 2.960 32.560 2.960
                 32.560 0.000 34.800 0.000 ;
        LAYER via3 ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal4 ;
        POLYGON  34.800 218.000 30.120 218.000 30.120 213.170 4.680 213.170 4.680 218.000
                 0.000 218.000 0.000 0.000 2.240 0.000 2.240 2.960 32.560 2.960
                 32.560 0.000 34.800 0.000 ;
        LAYER via4 ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal5 ;
        POLYGON  34.800 218.000 30.340 218.000 30.340 212.950 4.460 212.950 4.460 218.000
                 0.000 218.000 0.000 0.000 2.020 0.000 2.020 3.180 32.780 3.180
                 32.780 0.000 34.800 0.000 ;
        LAYER via5 ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal6 ;
        POLYGON  34.800 218.000 30.340 218.000 30.340 212.950 4.460 212.950 4.460 218.000
                 0.000 218.000 0.000 0.000 2.020 0.000 2.020 3.180 32.780 3.180
                 32.780 0.000 34.800 0.000 ;
        LAYER via6 ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal7 ;
        POLYGON  34.800 218.000 30.340 218.000 30.340 212.950 4.460 212.950 4.460 218.000
                 0.000 218.000 0.000 0.000 2.020 0.000 2.020 3.180 32.780 3.180
                 32.780 0.000 34.800 0.000 ;
        LAYER via7 ;
        RECT  2.520 0.000 32.280 2.680 ;
        RECT  4.960 213.450 29.840 218.000 ;
        LAYER metal8 ;
        POLYGON  34.800 218.000 30.340 218.000 30.340 212.950 4.460 212.950 4.460 218.000
                 0.000 218.000 0.000 0.000 2.020 0.000 2.020 3.180 32.780 3.180
                 32.780 0.000 34.800 0.000 ;
    END
END ULSCI0CUTHA

MACRO ULSCI0CUTHB
    CLASS PAD ;
    FOREIGN ULSCI0CUTHB 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 60.000 BY 152.000 ;
    SYMMETRY x y r90 ;
    SITE iocore_b ;
    PIN O
        DIRECTION INOUT ;
        PORT
        LAYER metal8 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal7 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal6 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal5 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal4 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal3 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal2 ;
        RECT  31.480 147.050 56.360 151.600 ;
        LAYER metal1 ;
        RECT  31.480 147.050 56.360 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal7 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal6 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal5 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal4 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal3 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal2 ;
        RECT  3.640 147.050 28.520 151.600 ;
        LAYER metal1 ;
        RECT  3.640 147.050 28.520 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal7 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal6 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal5 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal4 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal3 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal2 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal1 ;
        RECT  1.860 0.000 58.140 2.680 ;
        END
    END O
    PIN VCC12ANA
        DIRECTION INPUT ;
    END VCC12ANA
    PIN GNDANA
        DIRECTION INPUT ;
    END GNDANA
    OBS
        LAYER metal1 ;
        POLYGON  60.000 151.600 56.620 151.600 56.620 146.790 31.220 146.790
                 31.220 151.600 28.780 151.600 28.780 146.790 3.380 146.790 3.380 151.600
                 0.000 151.600 0.000 0.000 1.600 0.000 1.600 2.940 58.400 2.940
                 58.400 0.000 60.000 0.000 ;
        LAYER via ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal2 ;
        POLYGON  60.000 151.600 56.640 151.600 56.640 146.770 31.200 146.770
                 31.200 151.600 28.800 151.600 28.800 146.770 3.360 146.770 3.360 151.600
                 0.000 151.600 0.000 0.000 1.580 0.000 1.580 2.960 58.420 2.960
                 58.420 0.000 60.000 0.000 ;
        LAYER via2 ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal3 ;
        POLYGON  60.000 151.600 56.640 151.600 56.640 146.770 31.200 146.770
                 31.200 151.600 28.800 151.600 28.800 146.770 3.360 146.770 3.360 151.600
                 0.000 151.600 0.000 0.000 1.580 0.000 1.580 2.960 58.420 2.960
                 58.420 0.000 60.000 0.000 ;
        LAYER via3 ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal4 ;
        POLYGON  60.000 151.600 56.640 151.600 56.640 146.770 31.200 146.770
                 31.200 151.600 28.800 151.600 28.800 146.770 3.360 146.770 3.360 151.600
                 0.000 151.600 0.000 0.000 1.580 0.000 1.580 2.960 58.420 2.960
                 58.420 0.000 60.000 0.000 ;
        LAYER via4 ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal5 ;
        POLYGON  60.000 151.600 56.860 151.600 56.860 146.550 30.980 146.550
                 30.980 151.600 29.020 151.600 29.020 146.550 3.140 146.550 3.140 151.600
                 0.000 151.600 0.000 0.000 1.360 0.000 1.360 3.180 58.640 3.180
                 58.640 0.000 60.000 0.000 ;
        LAYER via5 ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal6 ;
        POLYGON  60.000 151.600 56.860 151.600 56.860 146.550 30.980 146.550
                 30.980 151.600 29.020 151.600 29.020 146.550 3.140 146.550 3.140 151.600
                 0.000 151.600 0.000 0.000 1.360 0.000 1.360 3.180 58.640 3.180
                 58.640 0.000 60.000 0.000 ;
        LAYER via6 ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal7 ;
        POLYGON  60.000 151.600 56.860 151.600 56.860 146.550 30.980 146.550
                 30.980 151.600 29.020 151.600 29.020 146.550 3.140 146.550 3.140 151.600
                 0.000 151.600 0.000 0.000 1.360 0.000 1.360 3.180 58.640 3.180
                 58.640 0.000 60.000 0.000 ;
        LAYER via7 ;
        RECT  31.480 147.050 56.360 151.600 ;
        RECT  3.640 147.050 28.520 151.600 ;
        RECT  1.860 0.000 58.140 2.680 ;
        LAYER metal8 ;
        POLYGON  60.000 151.600 56.860 151.600 56.860 146.550 30.980 146.550
                 30.980 151.600 29.020 151.600 29.020 146.550 3.140 146.550 3.140 151.600
                 0.000 151.600 0.000 0.000 1.360 0.000 1.360 3.180 58.640 3.180
                 58.640 0.000 60.000 0.000 ;
    END
END ULSCI0CUTHB

MACRO VCC12ACUTHA
    CLASS PAD ;
    FOREIGN VCC12ACUTHA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.800 BY 218.400 ;
    SYMMETRY x y r90 ;
    SITE iocore_a ;
    PIN VCC12ANA
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal7 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal6 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal5 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal4 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal3 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal2 ;
        RECT  22.080 213.450 38.280 218.000 ;
        LAYER metal1 ;
        RECT  22.080 213.450 38.280 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal7 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal6 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal5 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal4 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal3 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal2 ;
        RECT  2.520 213.450 18.720 218.000 ;
        LAYER metal1 ;
        RECT  2.520 213.450 18.720 218.000 ;
        END
        PORT
        LAYER metal8 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal7 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal6 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal5 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal4 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal3 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal2 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal1 ;
        RECT  2.000 0.000 38.800 3.480 ;
        END
    END VCC12ANA
    OBS
        LAYER metal1 ;
        POLYGON  40.800 218.000 38.540 218.000 38.540 213.190 21.820 213.190
                 21.820 218.000 18.980 218.000 18.980 213.190 2.260 213.190 2.260 218.000
                 0.000 218.000 0.000 0.000 1.740 0.000 1.740 3.740 39.060 3.740
                 39.060 0.000 40.800 0.000 ;
        LAYER via ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal2 ;
        POLYGON  40.800 218.000 38.560 218.000 38.560 213.170 21.800 213.170
                 21.800 218.000 19.000 218.000 19.000 213.170 2.240 213.170 2.240 218.000
                 0.000 218.000 0.000 0.000 1.720 0.000 1.720 3.760 39.080 3.760
                 39.080 0.000 40.800 0.000 ;
        LAYER via2 ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal3 ;
        POLYGON  40.800 218.000 38.560 218.000 38.560 213.170 21.800 213.170
                 21.800 218.000 19.000 218.000 19.000 213.170 2.240 213.170 2.240 218.000
                 0.000 218.000 0.000 0.000 1.720 0.000 1.720 3.760 39.080 3.760
                 39.080 0.000 40.800 0.000 ;
        LAYER via3 ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal4 ;
        POLYGON  40.800 218.000 38.560 218.000 38.560 213.170 21.800 213.170
                 21.800 218.000 19.000 218.000 19.000 213.170 2.240 213.170 2.240 218.000
                 0.000 218.000 0.000 0.000 1.720 0.000 1.720 3.760 39.080 3.760
                 39.080 0.000 40.800 0.000 ;
        LAYER via4 ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal5 ;
        POLYGON  40.800 218.000 38.780 218.000 38.780 212.950 21.580 212.950
                 21.580 218.000 19.220 218.000 19.220 212.950 2.020 212.950 2.020 218.000
                 0.000 218.000 0.000 0.000 1.500 0.000 1.500 3.980 39.300 3.980
                 39.300 0.000 40.800 0.000 ;
        LAYER via5 ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal6 ;
        POLYGON  40.800 218.000 38.780 218.000 38.780 212.950 21.580 212.950
                 21.580 218.000 19.220 218.000 19.220 212.950 2.020 212.950 2.020 218.000
                 0.000 218.000 0.000 0.000 1.500 0.000 1.500 3.980 39.300 3.980
                 39.300 0.000 40.800 0.000 ;
        LAYER via6 ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal7 ;
        POLYGON  40.800 218.000 38.780 218.000 38.780 212.950 21.580 212.950
                 21.580 218.000 19.220 218.000 19.220 212.950 2.020 212.950 2.020 218.000
                 0.000 218.000 0.000 0.000 1.500 0.000 1.500 3.980 39.300 3.980
                 39.300 0.000 40.800 0.000 ;
        LAYER via7 ;
        RECT  22.080 213.450 38.280 218.000 ;
        RECT  2.520 213.450 18.720 218.000 ;
        RECT  2.000 0.000 38.800 3.480 ;
        LAYER metal8 ;
        POLYGON  40.800 218.000 38.780 218.000 38.780 212.950 21.580 212.950
                 21.580 218.000 19.220 218.000 19.220 212.950 2.020 212.950 2.020 218.000
                 0.000 218.000 0.000 0.000 1.500 0.000 1.500 3.980 39.300 3.980
                 39.300 0.000 40.800 0.000 ;
    END
END VCC12ACUTHA

MACRO VCC12ACUTHB
    CLASS PAD ;
    FOREIGN VCC12ACUTHB 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.000 BY 152.000 ;
    SYMMETRY x y r90 ;
    SITE iocore_b ;
    PIN VCC12ANA
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal8 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal7 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal6 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal5 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal4 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal3 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal2 ;
        RECT  32.680 147.050 57.160 151.600 ;
        LAYER metal1 ;
        RECT  32.680 147.050 57.160 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal7 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal6 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal5 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal4 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal3 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal2 ;
        RECT  4.840 147.050 29.320 151.600 ;
        LAYER metal1 ;
        RECT  4.840 147.050 29.320 151.600 ;
        END
        PORT
        LAYER metal8 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal7 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal6 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal5 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal4 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal3 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal2 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal1 ;
        RECT  2.860 0.000 59.140 3.480 ;
        END
    END VCC12ANA
    OBS
        LAYER metal1 ;
        POLYGON  62.000 151.600 57.420 151.600 57.420 146.790 32.420 146.790
                 32.420 151.600 29.580 151.600 29.580 146.790 4.580 146.790 4.580 151.600
                 0.000 151.600 0.000 0.000 2.600 0.000 2.600 3.740 59.400 3.740
                 59.400 0.000 62.000 0.000 ;
        LAYER via ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal2 ;
        POLYGON  62.000 151.600 57.440 151.600 57.440 146.770 32.400 146.770
                 32.400 151.600 29.600 151.600 29.600 146.770 4.560 146.770 4.560 151.600
                 0.000 151.600 0.000 0.000 2.580 0.000 2.580 3.760 59.420 3.760
                 59.420 0.000 62.000 0.000 ;
        LAYER via2 ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal3 ;
        POLYGON  62.000 151.600 57.440 151.600 57.440 146.770 32.400 146.770
                 32.400 151.600 29.600 151.600 29.600 146.770 4.560 146.770 4.560 151.600
                 0.000 151.600 0.000 0.000 2.580 0.000 2.580 3.760 59.420 3.760
                 59.420 0.000 62.000 0.000 ;
        LAYER via3 ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal4 ;
        POLYGON  62.000 151.600 57.440 151.600 57.440 146.770 32.400 146.770
                 32.400 151.600 29.600 151.600 29.600 146.770 4.560 146.770 4.560 151.600
                 0.000 151.600 0.000 0.000 2.580 0.000 2.580 3.760 59.420 3.760
                 59.420 0.000 62.000 0.000 ;
        LAYER via4 ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal5 ;
        POLYGON  62.000 151.600 57.660 151.600 57.660 146.550 32.180 146.550
                 32.180 151.600 29.820 151.600 29.820 146.550 4.340 146.550 4.340 151.600
                 0.000 151.600 0.000 0.000 2.360 0.000 2.360 3.980 59.640 3.980
                 59.640 0.000 62.000 0.000 ;
        LAYER via5 ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal6 ;
        POLYGON  62.000 151.600 57.660 151.600 57.660 146.550 32.180 146.550
                 32.180 151.600 29.820 151.600 29.820 146.550 4.340 146.550 4.340 151.600
                 0.000 151.600 0.000 0.000 2.360 0.000 2.360 3.980 59.640 3.980
                 59.640 0.000 62.000 0.000 ;
        LAYER via6 ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal7 ;
        POLYGON  62.000 151.600 57.660 151.600 57.660 146.550 32.180 146.550
                 32.180 151.600 29.820 151.600 29.820 146.550 4.340 146.550 4.340 151.600
                 0.000 151.600 0.000 0.000 2.360 0.000 2.360 3.980 59.640 3.980
                 59.640 0.000 62.000 0.000 ;
        LAYER via7 ;
        RECT  32.680 147.050 57.160 151.600 ;
        RECT  4.840 147.050 29.320 151.600 ;
        RECT  2.860 0.000 59.140 3.480 ;
        LAYER metal8 ;
        POLYGON  62.000 151.600 57.660 151.600 57.660 146.550 32.180 146.550
                 32.180 151.600 29.820 151.600 29.820 146.550 4.340 146.550 4.340 151.600
                 0.000 151.600 0.000 0.000 2.360 0.000 2.360 3.980 59.640 3.980
                 59.640 0.000 62.000 0.000 ;
    END
END VCC12ACUTHB



END LIBRARY
