VERSION 5.5 ;
NAMESCASESENSITIVE ON ;




LAYER metal1  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal1

LAYER metal2
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal2

LAYER metal3
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal3

LAYER metal4  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal4

LAYER metal5  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal5

LAYER metal6
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal6

LAYER metal7  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1.1 ;  
END metal7

LAYER metal8  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1.1 ;  
END metal8


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:18 CST 2005
#
#**********************************************************************




MACRO AN2B1CHD
  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.688401 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.125600 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.442703 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.557600 LAYER metal1 ;
   AntennaDiffArea                            0.492000 LAYER metal1 ;
  END O

END AN2B1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:24 CST 2005
#
#**********************************************************************




MACRO AN2B1EHD
  PIN B1
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.360214 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.142000 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.266662 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AN2B1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:29 CST 2005
#
#**********************************************************************




MACRO AN2B1HHD
  PIN B1
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.360214 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.142000 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.904762 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.489600 LAYER metal1 ;
   AntennaDiffArea                            0.760800 LAYER metal1 ;
  END O

END AN2B1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:34 CST 2005
#
#**********************************************************************




MACRO AN2B1KHD
  PIN B1
   AntennaPartialMetalArea                    0.140000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.016667 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.367200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008714 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.820000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AN2B1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:39 CST 2005
#
#**********************************************************************




MACRO AN2CHD
  PIN I1
   AntennaPartialMetalArea                    0.131200 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.988888 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.988889 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.355200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AN2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:45 CST 2005
#
#**********************************************************************




MACRO AN2EHD
  PIN I1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.102000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.862744 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.102000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.917647 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AN2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:50 CST 2005
#
#**********************************************************************




MACRO AN2HHD
  PIN I1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.194400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.909464 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.194400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.880657 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.580800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AN2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:57:55 CST 2005
#
#**********************************************************************




MACRO AN2KHD
  PIN I1
   AntennaPartialMetalArea                    0.172000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.765959 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.336883 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.136000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AN2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:01 CST 2005
#
#**********************************************************************




MACRO AN3B1CHD
  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.069600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.229885 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.111600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.838707 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.111600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.788528 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.355200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END AN3B1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:06 CST 2005
#
#**********************************************************************




MACRO AN3B1EHD
  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.122224 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.040542 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.009005 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AN3B1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:11 CST 2005
#
#**********************************************************************




MACRO AN3B1HHD
  PIN B1
   AntennaPartialMetalArea                    0.140000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.291667 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.211200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.852271 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.211200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.825756 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.545600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AN3B1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:16 CST 2005
#
#**********************************************************************




MACRO AN3B2BHD
  PIN B1
   AntennaPartialMetalArea                    0.229600 LAYER metal1 ;
   AntennaGateArea                            0.162000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.202466 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.162000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.202467 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.122800 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.244444 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.682400 LAYER metal1 ;
   AntennaDiffArea                            0.682500 LAYER metal1 ;
  END O

END AN3B2BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:21 CST 2005
#
#**********************************************************************




MACRO AN3B2EHD
  PIN B1
   AntennaPartialMetalArea                    0.158800 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.505371 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.505380 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.123805 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AN3B2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:26 CST 2005
#
#**********************************************************************




MACRO AN3B2HHD
  PIN B1
   AntennaPartialMetalArea                    0.158800 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.849203 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.849209 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.881857 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.500800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AN3B2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:31 CST 2005
#
#**********************************************************************




MACRO AN3CHD
  PIN I1
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.349208 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.172800 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.071424 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.015872 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.355200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END AN3CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:36 CST 2005
#
#**********************************************************************




MACRO AN3EHD
  PIN I1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.487177 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.364105 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.160800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.256411 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.475200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AN3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:41 CST 2005
#
#**********************************************************************




MACRO AN3HHD
  PIN I1
   AntennaPartialMetalArea                    0.126400 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.112557 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.099566 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.146800 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.255408 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.475200 LAYER metal1 ;
   AntennaDiffArea                            0.883600 LAYER metal1 ;
  END O

END AN3HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:46 CST 2005
#
#**********************************************************************




MACRO AN4B1BHD
  PIN B1
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.138000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.281156 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.093600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.606841 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.172800 LAYER metal1 ;
   AntennaGateArea                            0.093600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.307696 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.093600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.247861 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.503600 LAYER metal1 ;
   AntennaDiffArea                            0.444000 LAYER metal1 ;
  END O

END AN4B1BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:52 CST 2005
#
#**********************************************************************




MACRO AN4B1EHD
  PIN B1
   AntennaPartialMetalArea                    0.816000 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.428569 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.323809 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.172800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.157139 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.123805 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.654000 LAYER metal1 ;
   AntennaDiffArea                            0.960000 LAYER metal1 ;
  END O

END AN4B1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:58:59 CST 2005
#
#**********************************************************************




MACRO AN4B1HHD
  PIN B1
   AntennaPartialMetalArea                    1.502400 LAYER metal1 ;
   AntennaGateArea                            0.691200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.552379 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.120000 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.112549 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.172800 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.961035 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.930740 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.504000 LAYER metal1 ;
   AntennaDiffArea                            1.808000 LAYER metal1 ;
  END O

END AN4B1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:08 CST 2005
#
#**********************************************************************




MACRO AN4CHD
  PIN I1
   AntennaPartialMetalArea                    0.131200 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.892469 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.892473 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.131200 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.892469 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.074400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.892477 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.408000 LAYER metal1 ;
   AntennaDiffArea                            0.926400 LAYER metal1 ;
  END O

END AN4CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:15 CST 2005
#
#**********************************************************************




MACRO AN4EHD
  PIN I1
   AntennaPartialMetalArea                    0.168000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.553330 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.553333 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.613337 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.156000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.753330 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.436000 LAYER metal1 ;
   AntennaDiffArea                            0.822400 LAYER metal1 ;
  END O

END AN4EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:20 CST 2005
#
#**********************************************************************




MACRO AN4HHD
  PIN I1
   AntennaPartialMetalArea                    0.172000 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.900902 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.027029 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.900904 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.156000 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.995492 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.244000 LAYER metal1 ;
   AntennaDiffArea                            1.644800 LAYER metal1 ;
  END O

END AN4HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:25 CST 2005
#
#**********************************************************************




MACRO ANTHD
  PIN A
   AntennaPartialMetalArea                    0.297600 LAYER metal1 ;
   AntennaDiffArea                            0.129600 LAYER metal1 ;
  END A

END ANTHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:36 CST 2005
#
#**********************************************************************




MACRO AO112CHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.191923 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.419196 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.983337 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.983333 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.355200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AO112CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:41 CST 2005
#
#**********************************************************************




MACRO AO112EHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.412126 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.383082 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911647 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911645 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AO112EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:46 CST 2005
#
#**********************************************************************




MACRO AO112HHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.412126 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.383082 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.866668 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.866663 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AO112HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:51 CST 2005
#
#**********************************************************************




MACRO AO112KHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.139200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287354 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.280952 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785181 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785182 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.179200 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AO112KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 20:59:56 CST 2005
#
#**********************************************************************




MACRO AO12CHD
  PIN A1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.793937 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.198063 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.164247 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.387200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AO12CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:00 CST 2005
#
#**********************************************************************




MACRO AO12EHD
  PIN A1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.048893 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.905978 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.933337 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AO12EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:05 CST 2005
#
#**********************************************************************




MACRO AO12HHD
  PIN A1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.102223 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783684 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758863 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.482000 LAYER metal1 ;
   AntennaDiffArea                            0.832000 LAYER metal1 ;
  END O

END AO12HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:10 CST 2005
#
#**********************************************************************




MACRO AO12KHD
  PIN A1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.995837 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783684 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758865 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.191200 LAYER metal1 ;
   AntennaDiffArea                            1.584000 LAYER metal1 ;
  END O

END AO12KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:16 CST 2005
#
#**********************************************************************




MACRO AO13CHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.136800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.362572 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.912701 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793646 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.793648 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.355200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AO13CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:20 CST 2005
#
#**********************************************************************




MACRO AO13EHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.151200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.105817 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AO13EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:25 CST 2005
#
#**********************************************************************




MACRO AO13HHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.151200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.105817 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AO13HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:30 CST 2005
#
#**********************************************************************




MACRO AO13KHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833333 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.179200 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AO13KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:35 CST 2005
#
#**********************************************************************




MACRO AO2222BHD
  PIN A1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.083337 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.213337 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.653337 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.746670 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.543333 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.066663 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.586670 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.586670 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.678000 LAYER metal1 ;
   AntennaDiffArea                            0.431200 LAYER metal1 ;
  END O

END AO2222BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:39 CST 2005
#
#**********************************************************************




MACRO AO2222CHD
  PIN A1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.842262 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.958337 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.458334 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.541667 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.377980 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755950 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.416667 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.416667 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.682000 LAYER metal1 ;
   AntennaDiffArea                            0.578200 LAYER metal1 ;
  END O

END AO2222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:44 CST 2005
#
#**********************************************************************




MACRO AO2222EHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.974076 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.113724 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740737 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792589 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740743 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.999997 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740739 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740737 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.998400 LAYER metal1 ;
   AntennaDiffArea                            0.892000 LAYER metal1 ;
  END O

END AO2222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:49 CST 2005
#
#**********************************************************************




MACRO AO2222HHD
  PIN A1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932621 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.113724 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709218 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758864 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.907797 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709217 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709222 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    1.523200 LAYER metal1 ;
   AntennaDiffArea                            1.581600 LAYER metal1 ;
  END O

END AO2222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:54 CST 2005
#
#**********************************************************************




MACRO AO222CHD
  PIN A1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.967588 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.126400 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.967589 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.226847 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.032409 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.097218 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.967589 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.299200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AO222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:00:59 CST 2005
#
#**********************************************************************




MACRO AO222EHD
  PIN A1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008333 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008330 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066663 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.891667 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.170400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.070421 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833337 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.475200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AO222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:04 CST 2005
#
#**********************************************************************




MACRO AO222HHD
  PIN A1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.894116 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839220 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.000005 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839218 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976467 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784314 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.519600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AO222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:09 CST 2005
#
#**********************************************************************




MACRO AO222KHD
  PIN A1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.894116 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839220 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.000005 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839218 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976467 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784314 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.999600 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AO222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:14 CST 2005
#
#**********************************************************************




MACRO AO22CHD
  PIN A1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.538687 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.505954 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.288687 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.288690 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.299200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AO22CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:18 CST 2005
#
#**********************************************************************




MACRO AO22EHD
  PIN A1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.896297 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.875923 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.896294 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740737 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.475200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AO22EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:23 CST 2005
#
#**********************************************************************




MACRO AO22HHD
  PIN A1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.808507 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758861 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.858153 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709222 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.520000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AO22HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:28 CST 2005
#
#**********************************************************************




MACRO AO22KHD
  PIN A1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.808514 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758868 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.858153 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709222 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.000000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AO22KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:32 CST 2005
#
#**********************************************************************




MACRO AOI112BHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.412126 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.383082 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911647 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911646 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.324000 LAYER metal1 ;
   AntennaDiffArea                            0.640000 LAYER metal1 ;
  END O

END AOI112BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:37 CST 2005
#
#**********************************************************************




MACRO AOI112EHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.191923 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.419196 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.983337 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.983337 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AOI112EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:41 CST 2005
#
#**********************************************************************




MACRO AOI112HHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.159209 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.383082 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911647 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911646 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.545600 LAYER metal1 ;
   AntennaDiffArea                            0.827200 LAYER metal1 ;
  END O

END AOI112HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:46 CST 2005
#
#**********************************************************************




MACRO AOI112KHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.159209 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.383082 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911647 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.911646 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.371200 LAYER metal1 ;
   AntennaDiffArea                            1.654400 LAYER metal1 ;
  END O

END AOI112KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:50 CST 2005
#
#**********************************************************************




MACRO AOI12CHD
  PIN A1
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.240433 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783686 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.126400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783686 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.244000 LAYER metal1 ;
   AntennaDiffArea                            0.873200 LAYER metal1 ;
  END O

END AOI12CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:01:55 CST 2005
#
#**********************************************************************




MACRO AOI12EHD
  PIN A1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.122400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.013072 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.343439 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.308085 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.505600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AOI12EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:00 CST 2005
#
#**********************************************************************




MACRO AOI12HHD
  PIN A1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.173520 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783684 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758865 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.577600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AOI12HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:05 CST 2005
#
#**********************************************************************




MACRO AOI12KHD
  PIN A1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.142224 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783684 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758865 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.259200 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AOI12KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:10 CST 2005
#
#**********************************************************************




MACRO AOI13BHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.133200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.399397 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.114400 LAYER metal1 ;
   AntennaDiffArea                            0.690600 LAYER metal1 ;
  END O

END AOI13BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:15 CST 2005
#
#**********************************************************************




MACRO AOI13EHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066662 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.467200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AOI13EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:20 CST 2005
#
#**********************************************************************




MACRO AOI13HHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.139200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287354 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.566400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AOI13HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:25 CST 2005
#
#**********************************************************************




MACRO AOI13KHD
  PIN A1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.139200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287354 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.815598 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709216 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709220 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.208000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AOI13KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:30 CST 2005
#
#**********************************************************************




MACRO AOI2222CHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.556414 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.656408 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.225642 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.297433 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.110259 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.461538 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.174358 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.174358 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.312400 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END AOI2222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:35 CST 2005
#
#**********************************************************************




MACRO AOI2222EHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.113724 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709222 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758867 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.957452 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758862 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758862 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.299200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AOI2222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:40 CST 2005
#
#**********************************************************************




MACRO AOI2222HHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.113724 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758867 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.957452 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758862 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758862 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.520000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AOI2222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:45 CST 2005
#
#**********************************************************************




MACRO AOI2222KHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.974076 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.113724 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740746 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792597 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740743 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.999997 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740739 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740737 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.936000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AOI2222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:50 CST 2005
#
#**********************************************************************




MACRO AOI222BHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.140559 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.887555 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.943780 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.943775 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.887550 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.887550 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.060000 LAYER metal1 ;
   AntennaDiffArea                            1.073200 LAYER metal1 ;
  END O

END AOI222BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:02:55 CST 2005
#
#**********************************************************************




MACRO AOI222EHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.979626 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.038886 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740746 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792597 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.075559 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.144800 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888886 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.475200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AOI222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:00 CST 2005
#
#**********************************************************************




MACRO AOI222HHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.994679 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758864 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.991565 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.178400 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.843882 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.520000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AOI222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:04 CST 2005
#
#**********************************************************************




MACRO AOI222KHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.007089 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758864 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.926833 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.178400 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.838416 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.936000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AOI222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:09 CST 2005
#
#**********************************************************************




MACRO AOI22BHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.130345 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.061402 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854700 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.914529 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.803200 LAYER metal1 ;
   AntennaDiffArea                            0.624000 LAYER metal1 ;
  END O

END AOI22BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:14 CST 2005
#
#**********************************************************************




MACRO AOI22EHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.979626 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.844447 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740746 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792597 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.475200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END AOI22EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:18 CST 2005
#
#**********************************************************************




MACRO AOI22HHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.960319 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758864 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.520000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END AOI22HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:24 CST 2005
#
#**********************************************************************




MACRO AOI22KHD
  PIN A1
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.858154 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758864 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.948000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END AOI22KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:29 CST 2005
#
#**********************************************************************




MACRO BHD1HD
  PIN H
   AntennaPartialMetalArea                    0.941600 LAYER metal1 ;
   AntennaGateArea                            1.579200 LAYER metal1 ;
   AntennaDiffArea                            0.217600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.588649 LAYER metal1 ; 
  END H

END BHD1HD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:33 CST 2005
#
#**********************************************************************




MACRO BUFBEHD
  PIN EB
   AntennaPartialMetalArea                    0.477600 LAYER metal1 ;
   AntennaGateArea                            0.352800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.418439 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.130400 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.075266 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaDiffArea                            0.672000 LAYER metal1 ;
  END O

END BUFBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:38 CST 2005
#
#**********************************************************************




MACRO BUFBHHD
  PIN EB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.401964 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.504660 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.532000 LAYER metal1 ;
   AntennaDiffArea                            0.672000 LAYER metal1 ;
  END O

END BUFBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:42 CST 2005
#
#**********************************************************************




MACRO BUFBIHD
  PIN EB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.401964 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.504660 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.708000 LAYER metal1 ;
   AntennaDiffArea                            1.154400 LAYER metal1 ;
  END O

END BUFBIHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:47 CST 2005
#
#**********************************************************************




MACRO BUFBKHD
  PIN EB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.401964 LAYER metal1 ; 
  END EB

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.504660 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.765600 LAYER metal1 ;
   AntennaDiffArea                            1.408000 LAYER metal1 ;
  END O

END BUFBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:51 CST 2005
#
#**********************************************************************




MACRO BUFCHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.070800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.276836 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.367200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END BUFCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:03:56 CST 2005
#
#**********************************************************************




MACRO BUFCKEHD
  PIN I
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.782047 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.432000 LAYER metal1 ;
   AntennaDiffArea                            0.418200 LAYER metal1 ;
  END O

END BUFCKEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:01 CST 2005
#
#**********************************************************************




MACRO BUFCKGHD
  PIN I
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.084612 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.528000 LAYER metal1 ;
   AntennaDiffArea                            0.452000 LAYER metal1 ;
  END O

END BUFCKGHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:05 CST 2005
#
#**********************************************************************




MACRO BUFCKHHD
  PIN I
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.195600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.057263 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.536000 LAYER metal1 ;
   AntennaDiffArea                            0.556000 LAYER metal1 ;
  END O

END BUFCKHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:11 CST 2005
#
#**********************************************************************




MACRO BUFCKIHD
  PIN I
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.235200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.933671 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.740200 LAYER metal1 ;
   AntennaDiffArea                            0.955600 LAYER metal1 ;
  END O

END BUFCKIHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:16 CST 2005
#
#**********************************************************************




MACRO BUFCKJHD
  PIN I
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.280800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.460118 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.767200 LAYER metal1 ;
   AntennaDiffArea                            1.091200 LAYER metal1 ;
  END O

END BUFCKJHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:21 CST 2005
#
#**********************************************************************




MACRO BUFCKKHD
  PIN I
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.391200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.575661 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.132400 LAYER metal1 ;
   AntennaDiffArea                            1.100000 LAYER metal1 ;
  END O

END BUFCKKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:27 CST 2005
#
#**********************************************************************




MACRO BUFCKLHD
  PIN I
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.492000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.752849 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.764800 LAYER metal1 ;
   AntennaDiffArea                            1.504800 LAYER metal1 ;
  END O

END BUFCKLHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:32 CST 2005
#
#**********************************************************************




MACRO BUFCKMHD
  PIN I
   AntennaPartialMetalArea                    0.188800 LAYER metal1 ;
   AntennaGateArea                            0.590400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.551487 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.079200 LAYER metal1 ;
   AntennaDiffArea                            1.652000 LAYER metal1 ;
  END O

END BUFCKMHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:37 CST 2005
#
#**********************************************************************




MACRO BUFCKNHD
  PIN I
   AntennaPartialMetalArea                    0.190400 LAYER metal1 ;
   AntennaGateArea                            0.787200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.573680 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.969600 LAYER metal1 ;
   AntennaDiffArea                            2.204000 LAYER metal1 ;
  END O

END BUFCKNHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:42 CST 2005
#
#**********************************************************************




MACRO BUFCKQHD
  PIN I
   AntennaPartialMetalArea                    0.542400 LAYER metal1 ;
   AntennaGateArea                            1.260000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.333654 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   10.995600 LAYER metal1 ;
   AntennaDiffArea                            4.932000 LAYER metal1 ;
  END O

END BUFCKQHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:46 CST 2005
#
#**********************************************************************




MACRO BUFDHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.070800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.276836 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.367200 LAYER metal1 ;
   AntennaDiffArea                            0.510000 LAYER metal1 ;
  END O

END BUFDHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:51 CST 2005
#
#**********************************************************************




MACRO BUFEHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.205560 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.367200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END BUFEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:04:56 CST 2005
#
#**********************************************************************




MACRO BUFGHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.114000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.845619 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.434400 LAYER metal1 ;
   AntennaDiffArea                            0.600000 LAYER metal1 ;
  END O

END BUFGHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:01 CST 2005
#
#**********************************************************************




MACRO BUFHHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.134400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.565472 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.434400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END BUFHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:05 CST 2005
#
#**********************************************************************




MACRO BUFIHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.138531 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.745600 LAYER metal1 ;
   AntennaDiffArea                            1.165600 LAYER metal1 ;
  END O

END BUFIHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:10 CST 2005
#
#**********************************************************************




MACRO BUFJHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932624 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.699200 LAYER metal1 ;
   AntennaDiffArea                            1.401600 LAYER metal1 ;
  END O

END BUFJHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:15 CST 2005
#
#**********************************************************************




MACRO BUFKHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.301200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.580342 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.734400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END BUFKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:20 CST 2005
#
#**********************************************************************




MACRO BUFLHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.368400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.187840 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.024000 LAYER metal1 ;
   AntennaDiffArea                            2.143200 LAYER metal1 ;
  END O

END BUFLHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:25 CST 2005
#
#**********************************************************************




MACRO BUFMHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.444000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.985584 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.067200 LAYER metal1 ;
   AntennaDiffArea                            2.256000 LAYER metal1 ;
  END O

END BUFMHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:30 CST 2005
#
#**********************************************************************




MACRO BUFNHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.590400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.220868 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.096000 LAYER metal1 ;
   AntennaDiffArea                            3.008000 LAYER metal1 ;
  END O

END BUFNHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:35 CST 2005
#
#**********************************************************************




MACRO BUFQHD
  PIN I
   AntennaPartialMetalArea                    1.008000 LAYER metal1 ;
   AntennaGateArea                            1.488000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.310751 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   11.213200 LAYER metal1 ;
   AntennaDiffArea                            7.520000 LAYER metal1 ;
  END O

END BUFQHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:40 CST 2005
#
#**********************************************************************




MACRO BUFTEHD
  PIN E
   AntennaPartialMetalArea                    0.477600 LAYER metal1 ;
   AntennaGateArea                            0.271200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.481478 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.130400 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.075266 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.320000 LAYER metal1 ;
   AntennaDiffArea                            0.672000 LAYER metal1 ;
  END O

END BUFTEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:45 CST 2005
#
#**********************************************************************




MACRO BUFTHHD
  PIN E
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.240000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.635000 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.413750 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.536000 LAYER metal1 ;
   AntennaDiffArea                            0.672000 LAYER metal1 ;
  END O

END BUFTHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:50 CST 2005
#
#**********************************************************************




MACRO BUFTIHD
  PIN E
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.240000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.635000 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.343200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.413750 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.702400 LAYER metal1 ;
   AntennaDiffArea                            1.154400 LAYER metal1 ;
  END O

END BUFTIHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:54 CST 2005
#
#**********************************************************************




MACRO BUFTJHD
  PIN E
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.583334 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.354000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.357060 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.702400 LAYER metal1 ;
   AntennaDiffArea                            1.128000 LAYER metal1 ;
  END O

END BUFTJHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:05:59 CST 2005
#
#**********************************************************************




MACRO BUFTKHD
  PIN E
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.583334 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.354000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.377400 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.702400 LAYER metal1 ;
   AntennaDiffArea                            1.408000 LAYER metal1 ;
  END O

END BUFTKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:04 CST 2005
#
#**********************************************************************




MACRO CKLDHD
  PIN I
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.153504 LAYER metal1 ; 
  END I

END CKLDHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:09 CST 2005
#
#**********************************************************************




MACRO DBAHRBEHD
  PIN D
   AntennaPartialMetalArea                    0.163200 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.076581 LAYER metal1 ; 
  END D

  PIN GB
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END GB

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.446800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.135200 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976195 LAYER metal1 ; 
  END RB

END DBAHRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:15 CST 2005
#
#**********************************************************************




MACRO DBAHRBHHD
  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.033752 LAYER metal1 ; 
  END D

  PIN GB
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.603770 LAYER metal1 ; 
  END GB

  PIN Q
   AntennaPartialMetalArea                    0.332400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.392000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.130000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.063489 LAYER metal1 ; 
  END RB

END DBAHRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:19 CST 2005
#
#**********************************************************************




MACRO DBFRBEHD
  PIN CKB
   AntennaPartialMetalArea                    0.147600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609929 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.339200 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

END DBFRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:24 CST 2005
#
#**********************************************************************




MACRO DBFRBHHD
  PIN CKB
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609932 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.302000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.392400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

END DBFRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:29 CST 2005
#
#**********************************************************************




MACRO DBFRSBEHD
  PIN CKB
   AntennaPartialMetalArea                    0.138800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.613474 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.104170 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.411200 LAYER metal1 ;
   AntennaDiffArea                            0.575200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.165000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.268819 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.110800 LAYER metal1 ;
   AntennaGateArea                            0.153600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.057296 LAYER metal1 ; 
  END SB

END DBFRSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:35 CST 2005
#
#**********************************************************************




MACRO DBFRSBHHD
  PIN CKB
   AntennaPartialMetalArea                    0.138800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.133330 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.337600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.126000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.673204 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.138000 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.583333 LAYER metal1 ; 
  END SB

END DBFRSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:39 CST 2005
#
#**********************************************************************




MACRO DBZRBEHD
  PIN CKB
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.631202 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.344000 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END DBZRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:44 CST 2005
#
#**********************************************************************




MACRO DBZRBHHD
  PIN CKB
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.631202 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.302000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.392400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490433 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END DBZRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:49 CST 2005
#
#**********************************************************************




MACRO DBZRSBEHD
  PIN CKB
   AntennaPartialMetalArea                    0.110800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634750 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.944449 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.321600 LAYER metal1 ;
   AntennaDiffArea                            0.555200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.150000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.413975 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.153600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.057288 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.194000 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.463767 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.202381 LAYER metal1 ; 
  END TD

END DBZRSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:53 CST 2005
#
#**********************************************************************




MACRO DBZRSBHHD
  PIN CKB
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609931 LAYER metal1 ; 
  END CKB

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854699 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.337600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.126000 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.624184 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.122000 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.577269 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.670289 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.404761 LAYER metal1 ; 
  END TD

END DBZRSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:06:58 CST 2005
#
#**********************************************************************




MACRO DELAKHD
  PIN I
   AntennaPartialMetalArea                    0.228400 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.840579 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.120000 LAYER metal1 ;
   AntennaDiffArea                            1.584000 LAYER metal1 ;
  END O

END DELAKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:03 CST 2005
#
#**********************************************************************




MACRO DELBKHD
  PIN I
   AntennaPartialMetalArea                    0.228400 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.840579 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.120000 LAYER metal1 ;
   AntennaDiffArea                            1.584000 LAYER metal1 ;
  END O

END DELBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:08 CST 2005
#
#**********************************************************************




MACRO DELCKHD
  PIN I
   AntennaPartialMetalArea                    0.228400 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.840579 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.120000 LAYER metal1 ;
   AntennaDiffArea                            1.584000 LAYER metal1 ;
  END O

END DELCKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:12 CST 2005
#
#**********************************************************************




MACRO DELDKHD
  PIN I
   AntennaPartialMetalArea                    0.228400 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.840579 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.120000 LAYER metal1 ;
   AntennaDiffArea                            1.584000 LAYER metal1 ;
  END O

END DELDKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:17 CST 2005
#
#**********************************************************************




MACRO DFCLRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888886 LAYER metal1 ; 
  END D

  PIN LD
   AntennaPartialMetalArea                    0.780800 LAYER metal1 ;
   AntennaGateArea                            0.271200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.810254 LAYER metal1 ; 
  END LD

  PIN Q
   AntennaPartialMetalArea                    0.385600 LAYER metal1 ;
   AntennaDiffArea                            0.485200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.021372 LAYER metal1 ; 
  END RB

END DFCLRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:22 CST 2005
#
#**********************************************************************




MACRO DFCLRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888886 LAYER metal1 ; 
  END D

  PIN LD
   AntennaPartialMetalArea                    0.780800 LAYER metal1 ;
   AntennaGateArea                            0.271200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.810254 LAYER metal1 ; 
  END LD

  PIN Q
   AntennaPartialMetalArea                    0.293600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.382400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.021372 LAYER metal1 ; 
  END RB

END DFCLRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:27 CST 2005
#
#**********************************************************************




MACRO DFCRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.138800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.592204 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.616353 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.497200 LAYER metal1 ;
   AntennaDiffArea                            0.479600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.025158 LAYER metal1 ; 
  END RB

END DFCRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:32 CST 2005
#
#**********************************************************************




MACRO DFCRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.138800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.592204 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.616353 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.293600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.382400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.025158 LAYER metal1 ; 
  END RB

END DFCRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:37 CST 2005
#
#**********************************************************************




MACRO DFECHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.408890 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.292800 LAYER metal1 ;
   AntennaDiffArea                            0.302400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.278400 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END QB

END DFECHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:42 CST 2005
#
#**********************************************************************




MACRO DFEEHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.858157 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.326400 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

END DFEEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:47 CST 2005
#
#**********************************************************************




MACRO DFEHHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.858157 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.232000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.382400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

END DFEHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:52 CST 2005
#
#**********************************************************************




MACRO DFEKHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833337 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.792000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.792000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

END DFEKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:07:57 CST 2005
#
#**********************************************************************




MACRO DFERBCHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.142222 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.388800 LAYER metal1 ;
   AntennaDiffArea                            0.367600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.179400 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.838705 LAYER metal1 ; 
  END RB

END DFERBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:02 CST 2005
#
#**********************************************************************




MACRO DFERBEHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaDiffArea                            0.575200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.179400 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.416175 LAYER metal1 ; 
  END RB

END DFERBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:07 CST 2005
#
#**********************************************************************




MACRO DFERBHHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.243200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.363200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.179400 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.316935 LAYER metal1 ; 
  END RB

END DFERBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:12 CST 2005
#
#**********************************************************************




MACRO DFERBKHD
  PIN CK
   AntennaPartialMetalArea                    0.139600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.721636 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.792000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.792000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.152000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.481214 LAYER metal1 ; 
  END RB

END DFERBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:17 CST 2005
#
#**********************************************************************




MACRO DFERSBCHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.128892 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.268800 LAYER metal1 ;
   AntennaDiffArea                            0.367600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.205000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.091402 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.989740 LAYER metal1 ; 
  END SB

END DFERSBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:23 CST 2005
#
#**********************************************************************




MACRO DFERSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaDiffArea                            0.575200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.205000 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.471543 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.989740 LAYER metal1 ; 
  END SB

END DFERSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:28 CST 2005
#
#**********************************************************************




MACRO DFERSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.337600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.105600 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.717317 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.704549 LAYER metal1 ; 
  END SB

END DFERSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:33 CST 2005
#
#**********************************************************************




MACRO DFERSBKHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.721627 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.156400 LAYER metal1 ;
   AntennaGateArea                            0.126000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.755560 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.214800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.922718 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.123600 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.717318 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.601515 LAYER metal1 ; 
  END SB

END DFERSBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:37 CST 2005
#
#**********************************************************************




MACRO DFFCHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.128890 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.371200 LAYER metal1 ;
   AntennaDiffArea                            0.330400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END QB

END DFFCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:42 CST 2005
#
#**********************************************************************




MACRO DFFEHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570923 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.371200 LAYER metal1 ;
   AntennaDiffArea                            0.485200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

END DFFEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:47 CST 2005
#
#**********************************************************************




MACRO DFFHHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.393600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.332800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

END DFFHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:52 CST 2005
#
#**********************************************************************




MACRO DFFKHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.808000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.814400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

END DFFKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:08:57 CST 2005
#
#**********************************************************************




MACRO DFFRBCHD
  PIN CK
   AntennaPartialMetalArea                    0.147600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.177780 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.375600 LAYER metal1 ;
   AntennaDiffArea                            0.328600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

END DFFRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:01 CST 2005
#
#**********************************************************************




MACRO DFFRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.147600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609929 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.339200 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

END DFFRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:06 CST 2005
#
#**********************************************************************




MACRO DFFRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843967 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.302000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.392400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

END DFFRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:11 CST 2005
#
#**********************************************************************




MACRO DFFRBKHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709217 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.086400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.080000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

END DFFRBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:16 CST 2005
#
#**********************************************************************




MACRO DFFRSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634752 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.112497 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.253600 LAYER metal1 ;
   AntennaDiffArea                            0.575200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.205000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.268822 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.116400 LAYER metal1 ;
   AntennaGateArea                            0.153600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.088538 LAYER metal1 ; 
  END SB

END DFFRSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:21 CST 2005
#
#**********************************************************************




MACRO DFFRSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634752 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.112497 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.337600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.105600 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.638887 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.590909 LAYER metal1 ; 
  END SB

END DFFRSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:26 CST 2005
#
#**********************************************************************




MACRO DFFSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609932 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.364000 LAYER metal1 ;
   AntennaDiffArea                            0.580400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.300800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN SB
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.237600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.077440 LAYER metal1 ; 
  END SB

END DFFSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:30 CST 2005
#
#**********************************************************************




MACRO DFFSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609932 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.264000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.390400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN SB
   AntennaPartialMetalArea                    0.118000 LAYER metal1 ;
   AntennaGateArea                            0.319200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.174186 LAYER metal1 ; 
  END SB

END DFFSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:35 CST 2005
#
#**********************************************************************




MACRO DFTRBCHD
  PIN CK
   AntennaPartialMetalArea                    0.167600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.177778 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.036529 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.440000 LAYER metal1 ;
   AntennaDiffArea                            0.341200 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.258000 LAYER metal1 ;
   AntennaDiffArea                            0.446400 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

END DFTRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:40 CST 2005
#
#**********************************************************************




MACRO DFTRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.167600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.684394 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.276000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.214491 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.299200 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.400000 LAYER metal1 ;
   AntennaDiffArea                            0.736000 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

END DFTRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:46 CST 2005
#
#**********************************************************************




MACRO DFZCHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.128890 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.396800 LAYER metal1 ;
   AntennaDiffArea                            0.358400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END DFZCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:09:51 CST 2005
#
#**********************************************************************




MACRO DFZCLRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888886 LAYER metal1 ; 
  END D

  PIN LD
   AntennaPartialMetalArea                    0.707200 LAYER metal1 ;
   AntennaGateArea                            0.271200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.810260 LAYER metal1 ; 
  END LD

  PIN Q
   AntennaPartialMetalArea                    0.385600 LAYER metal1 ;
   AntennaDiffArea                            0.485200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854702 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.151200 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.440217 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.158000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.750000 LAYER metal1 ; 
  END TD

END DFZCLRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:02 CST 2005
#
#**********************************************************************




MACRO DFZCLRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888886 LAYER metal1 ; 
  END D

  PIN LD
   AntennaPartialMetalArea                    0.707200 LAYER metal1 ;
   AntennaGateArea                            0.271200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.810260 LAYER metal1 ; 
  END LD

  PIN Q
   AntennaPartialMetalArea                    0.293600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.382400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854702 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.151200 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.440217 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.158000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.750000 LAYER metal1 ; 
  END TD

END DFZCLRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:07 CST 2005
#
#**********************************************************************




MACRO DFZCRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.138800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.592204 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.390355 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.497200 LAYER metal1 ;
   AntennaDiffArea                            0.479600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267545 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.723000 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.595233 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.827385 LAYER metal1 ; 
  END TD

END DFZCRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:17 CST 2005
#
#**********************************************************************




MACRO DFZCRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.138800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.592204 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.390355 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.293600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.382400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267545 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.723000 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.595233 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.827385 LAYER metal1 ; 
  END TD

END DFZCRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:23 CST 2005
#
#**********************************************************************




MACRO DFZECHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.017780 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.280800 LAYER metal1 ;
   AntennaDiffArea                            0.330400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZECHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:28 CST 2005
#
#**********************************************************************




MACRO DFZEEHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609933 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.280800 LAYER metal1 ;
   AntennaDiffArea                            0.482400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZEEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:33 CST 2005
#
#**********************************************************************




MACRO DFZEHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.385600 LAYER metal1 ;
   AntennaDiffArea                            0.485200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.319200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END DFZEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:43 CST 2005
#
#**********************************************************************




MACRO DFZEHHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.546103 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.305600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.362400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZEHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:48 CST 2005
#
#**********************************************************************




MACRO DFZEKHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709217 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.882000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.948000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.459122 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZEKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:53 CST 2005
#
#**********************************************************************




MACRO DFZERBCHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.142222 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.388800 LAYER metal1 ;
   AntennaDiffArea                            0.367600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.179400 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.838705 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:10:58 CST 2005
#
#**********************************************************************




MACRO DFZERBEHD
  PIN CK
   AntennaPartialMetalArea                    0.136000 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.808506 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaDiffArea                            0.575200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.345172 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.421382 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:03 CST 2005
#
#**********************************************************************




MACRO DFZERBHHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.243200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.363200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.179400 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.316935 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:08 CST 2005
#
#**********************************************************************




MACRO DFZERBKHD
  PIN CK
   AntennaPartialMetalArea                    0.139600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.721636 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.152000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.481214 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.430822 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:14 CST 2005
#
#**********************************************************************




MACRO DFZERSBCHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.128892 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.268800 LAYER metal1 ;
   AntennaDiffArea                            0.367600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.205000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.091402 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.989740 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERSBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:18 CST 2005
#
#**********************************************************************




MACRO DFZERSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.285600 LAYER metal1 ;
   AntennaDiffArea                            0.575200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.205000 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.471543 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.989740 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:23 CST 2005
#
#**********************************************************************




MACRO DFZERSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634754 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.337600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.105600 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.717317 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.704549 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.477992 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:28 CST 2005
#
#**********************************************************************




MACRO DFZERSBKHD
  PIN CK
   AntennaPartialMetalArea                    0.127600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.721627 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273222 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.681162 LAYER metal1 ; 
  END EB

  PIN Q
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.123600 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.717318 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.601515 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.254400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.430822 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.404372 LAYER metal1 ; 
  END TD

END DFZERSBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:44 CST 2005
#
#**********************************************************************




MACRO DFZHHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.393600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.332800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END DFZHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:11:58 CST 2005
#
#**********************************************************************




MACRO DFZKHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.808000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.814400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END DFZKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:03 CST 2005
#
#**********************************************************************




MACRO DFZRBCHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.311110 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.281600 LAYER metal1 ;
   AntennaDiffArea                            0.367600 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.095239 LAYER metal1 ; 
  END TD

END DFZRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:08 CST 2005
#
#**********************************************************************




MACRO DFZRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.968083 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.344000 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721892 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END DFZRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:24 CST 2005
#
#**********************************************************************




MACRO DFZRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843967 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.302000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.392400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END DFZRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:34 CST 2005
#
#**********************************************************************




MACRO DFZRBKHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.086400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    1.080000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END DFZRBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:39 CST 2005
#
#**********************************************************************




MACRO DFZRSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.110800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634750 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.918799 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.321600 LAYER metal1 ;
   AntennaDiffArea                            0.555200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.259200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.160000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.413981 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.153600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.088537 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.507249 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.309521 LAYER metal1 ; 
  END TD

END DFZRSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:44 CST 2005
#
#**********************************************************************




MACRO DFZRSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634752 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854699 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.276800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.337600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.105600 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.638887 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.264000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.590909 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.670289 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.404761 LAYER metal1 ; 
  END TD

END DFZRSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:49 CST 2005
#
#**********************************************************************




MACRO DFZSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.116400 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609925 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854699 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.377600 LAYER metal1 ;
   AntennaDiffArea                            0.580400 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN SB
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.237600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158247 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.670289 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.404761 LAYER metal1 ; 
  END TD

END DFZSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:54 CST 2005
#
#**********************************************************************




MACRO DFZSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609932 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854699 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.264000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.390400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN SB
   AntennaPartialMetalArea                    0.118000 LAYER metal1 ;
   AntennaGateArea                            0.319200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.174186 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.670289 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.404761 LAYER metal1 ; 
  END TD

END DFZSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:12:59 CST 2005
#
#**********************************************************************




MACRO DFZTRBCHD
  PIN CK
   AntennaPartialMetalArea                    0.178800 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.271113 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.885849 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.344000 LAYER metal1 ;
   AntennaDiffArea                            0.302400 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.276000 LAYER metal1 ;
   AntennaDiffArea                            0.459000 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721889 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.136400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583336 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.041663 LAYER metal1 ; 
  END TD

END DFZTRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:04 CST 2005
#
#**********************************************************************




MACRO DFZTRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.178800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.684394 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.149600 LAYER metal1 ;
   AntennaGateArea                            0.276000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.214491 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.299200 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN QZ
   AntennaPartialMetalArea                    0.400000 LAYER metal1 ;
   AntennaDiffArea                            0.736000 LAYER metal1 ;
  END QZ

  PIN RB
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.721889 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.136400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583336 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.041663 LAYER metal1 ; 
  END TD

END DFZTRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:09 CST 2005
#
#**********************************************************************




MACRO DLAHCHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.688402 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.352800 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END QB

END DLAHCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:14 CST 2005
#
#**********************************************************************




MACRO DLAHEHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.139200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.347696 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.448800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

END DLAHEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:19 CST 2005
#
#**********************************************************************




MACRO DLAHHHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783690 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.603770 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.326800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.460000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

END DLAHHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:24 CST 2005
#
#**********************************************************************




MACRO DLAHRBCHD
  PIN D
   AntennaPartialMetalArea                    0.163200 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.076581 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.091200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.710530 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.352800 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.135200 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976195 LAYER metal1 ; 
  END RB

END DLAHRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:29 CST 2005
#
#**********************************************************************




MACRO DLAHRBEHD
  PIN D
   AntennaPartialMetalArea                    0.163200 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008441 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.446800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.135200 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976195 LAYER metal1 ; 
  END RB

END DLAHRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:34 CST 2005
#
#**********************************************************************




MACRO DLAHRBHHD
  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.912699 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.603770 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.332400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN QB
   AntennaPartialMetalArea                    0.392000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END QB

  PIN RB
   AntennaPartialMetalArea                    0.130000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.063489 LAYER metal1 ; 
  END RB

END DLAHRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:39 CST 2005
#
#**********************************************************************




MACRO FA1DHD
  PIN A
   AntennaPartialMetalArea                    1.192000 LAYER metal1 ;
   AntennaGateArea                            0.612000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.143628 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.157600 LAYER metal1 ;
   AntennaGateArea                            0.650400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.020322 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    1.344400 LAYER metal1 ;
   AntennaGateArea                            0.445200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.767024 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    0.283200 LAYER metal1 ;
   AntennaDiffArea                            0.578000 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.363200 LAYER metal1 ;
   AntennaDiffArea                            0.503200 LAYER metal1 ;
  END S

END FA1DHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:44 CST 2005
#
#**********************************************************************




MACRO FA1EHD
  PIN A
   AntennaPartialMetalArea                    0.494400 LAYER metal1 ;
   AntennaGateArea                            0.468000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.517950 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.509600 LAYER metal1 ;
   AntennaGateArea                            0.535200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.143373 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    2.096200 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.948710 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    0.387200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.377200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END S

END FA1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:49 CST 2005
#
#**********************************************************************




MACRO FA1HHD
  PIN A
   AntennaPartialMetalArea                    0.542800 LAYER metal1 ;
   AntennaGateArea                            0.468000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.466671 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.550000 LAYER metal1 ;
   AntennaGateArea                            0.564000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.726983 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    2.104800 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.595204 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    0.520000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.568000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END S

END FA1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:53 CST 2005
#
#**********************************************************************




MACRO FA1KHD
  PIN A
   AntennaPartialMetalArea                    0.542800 LAYER metal1 ;
   AntennaGateArea                            0.583200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.381643 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.517200 LAYER metal1 ;
   AntennaGateArea                            0.748800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.966185 LAYER metal1 ; 
  END B

  PIN CI
   AntennaPartialMetalArea                    2.108800 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.418519 LAYER metal1 ; 
  END CI

  PIN CO
   AntennaPartialMetalArea                    0.952000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END CO

  PIN S
   AntennaPartialMetalArea                    0.936000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END S

END FA1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:13:58 CST 2005
#
#**********************************************************************




MACRO GCBETCHD
  PIN CKB
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.122400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.385617 LAYER metal1 ; 
  END CKB

  PIN E
   AntennaPartialMetalArea                    0.220000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.191663 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.592800 LAYER metal1 ;
   AntennaDiffArea                            0.934400 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.144400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.915660 LAYER metal1 ; 
  END TE

END GCBETCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:03 CST 2005
#
#**********************************************************************




MACRO GCBETEHD
  PIN CKB
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.122400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.385617 LAYER metal1 ; 
  END CKB

  PIN E
   AntennaPartialMetalArea                    0.220000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.191663 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.308800 LAYER metal1 ;
   AntennaDiffArea                            0.489600 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.144400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.915660 LAYER metal1 ; 
  END TE

END GCBETEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:08 CST 2005
#
#**********************************************************************




MACRO GCBETHHD
  PIN CKB
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.122400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.385617 LAYER metal1 ; 
  END CKB

  PIN E
   AntennaPartialMetalArea                    0.220000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.191663 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.370400 LAYER metal1 ;
   AntennaDiffArea                            0.576000 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.161200 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.933733 LAYER metal1 ; 
  END TE

END GCBETHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:13 CST 2005
#
#**********************************************************************




MACRO GCBETKHD
  PIN CKB
   AntennaPartialMetalArea                    0.133600 LAYER metal1 ;
   AntennaGateArea                            0.122400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.385617 LAYER metal1 ; 
  END CKB

  PIN E
   AntennaPartialMetalArea                    0.220000 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.191663 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.692000 LAYER metal1 ;
   AntennaDiffArea                            1.152000 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.161200 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.933733 LAYER metal1 ; 
  END TE

END GCBETKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:18 CST 2005
#
#**********************************************************************




MACRO GCKETCHD
  PIN CK
   AntennaPartialMetalArea                    0.552000 LAYER metal1 ;
   AntennaGateArea                            0.321600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.581702 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.308337 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.319600 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.128400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.803212 LAYER metal1 ; 
  END TE

END GCKETCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:23 CST 2005
#
#**********************************************************************




MACRO GCKETEHD
  PIN CK
   AntennaPartialMetalArea                    0.552000 LAYER metal1 ;
   AntennaGateArea                            0.321600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.581702 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.308337 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.321200 LAYER metal1 ;
   AntennaDiffArea                            0.489600 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.128400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.803212 LAYER metal1 ; 
  END TE

END GCKETEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:28 CST 2005
#
#**********************************************************************




MACRO GCKETHHD
  PIN CK
   AntennaPartialMetalArea                    0.552000 LAYER metal1 ;
   AntennaGateArea                            0.321600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.581702 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.308337 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    0.745600 LAYER metal1 ;
   AntennaDiffArea                            0.979200 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.128400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.803212 LAYER metal1 ; 
  END TE

END GCKETHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:14:32 CST 2005
#
#**********************************************************************




MACRO GCKETKHD
  PIN CK
   AntennaPartialMetalArea                    0.552000 LAYER metal1 ;
   AntennaGateArea                            0.321600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.581702 LAYER metal1 ; 
  END CK

  PIN E
   AntennaPartialMetalArea                    0.231200 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.308337 LAYER metal1 ; 
  END E

  PIN Q
   AntennaPartialMetalArea                    1.123200 LAYER metal1 ;
   AntennaDiffArea                            1.555200 LAYER metal1 ;
  END Q

  PIN TE
   AntennaPartialMetalArea                    0.128400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.803212 LAYER metal1 ; 
  END TE

END GCKETKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:17 CST 2005
#
#**********************************************************************




MACRO HA1CHD
  PIN A
   AntennaPartialMetalArea                    0.115600 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.412935 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.008000 LAYER metal1 ;
   AntennaGateArea                            0.208800 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.031744 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.473600 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.369200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END S

END HA1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:21 CST 2005
#
#**********************************************************************




MACRO HA1EHD
  PIN A
   AntennaPartialMetalArea                    0.115600 LAYER metal1 ;
   AntennaGateArea                            0.230400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.913194 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.022400 LAYER metal1 ;
   AntennaGateArea                            0.283200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.757581 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.354400 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.371200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END S

END HA1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:26 CST 2005
#
#**********************************************************************




MACRO HA1HHD
  PIN A
   AntennaPartialMetalArea                    0.642800 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.651109 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.236000 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.366672 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.360000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END S

END HA1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:31 CST 2005
#
#**********************************************************************




MACRO HA1KHD
  PIN A
   AntennaPartialMetalArea                    0.719600 LAYER metal1 ;
   AntennaGateArea                            0.388800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.259467 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    1.300000 LAYER metal1 ;
   AntennaGateArea                            0.410400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.546299 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.614400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END C

  PIN S
   AntennaPartialMetalArea                    0.732800 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END S

END HA1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:35 CST 2005
#
#**********************************************************************




MACRO INVCHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.135600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.410030 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.351200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END INVCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:40 CST 2005
#
#**********************************************************************




MACRO INVCKDHD
  PIN I
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.129600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.790123 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.382800 LAYER metal1 ;
   AntennaDiffArea                            0.496800 LAYER metal1 ;
  END O

END INVCKDHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:45 CST 2005
#
#**********************************************************************




MACRO INVCKGHD
  PIN I
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.246000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.668290 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.500000 LAYER metal1 ;
   AntennaDiffArea                            0.495000 LAYER metal1 ;
  END O

END INVCKGHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:50 CST 2005
#
#**********************************************************************




MACRO INVCKHHD
  PIN I
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.328800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.508518 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.652000 LAYER metal1 ;
   AntennaDiffArea                            0.548000 LAYER metal1 ;
  END O

END INVCKHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:55 CST 2005
#
#**********************************************************************




MACRO INVCKIHD
  PIN I
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.405600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.806706 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.864000 LAYER metal1 ;
   AntennaDiffArea                            0.884000 LAYER metal1 ;
  END O

END INVCKIHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:15:59 CST 2005
#
#**********************************************************************




MACRO INVCKJHD
  PIN I
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.488400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.809994 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.024800 LAYER metal1 ;
   AntennaDiffArea                            1.045000 LAYER metal1 ;
  END O

END INVCKJHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:04 CST 2005
#
#**********************************************************************




MACRO INVCKKHD
  PIN I
   AntennaPartialMetalArea                    0.140800 LAYER metal1 ;
   AntennaGateArea                            0.652800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.598044 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.316400 LAYER metal1 ;
   AntennaDiffArea                            1.088000 LAYER metal1 ;
  END O

END INVCKKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:09 CST 2005
#
#**********************************************************************




MACRO INVCKLHD
  PIN I
   AntennaPartialMetalArea                    0.226000 LAYER metal1 ;
   AntennaGateArea                            0.819600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.601756 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.168200 LAYER metal1 ;
   AntennaDiffArea                            1.557800 LAYER metal1 ;
  END O

END INVCKLHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:15 CST 2005
#
#**********************************************************************




MACRO INVCKMHD
  PIN I
   AntennaPartialMetalArea                    0.256000 LAYER metal1 ;
   AntennaGateArea                            0.982800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.628000 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.402400 LAYER metal1 ;
   AntennaDiffArea                            1.639000 LAYER metal1 ;
  END O

END INVCKMHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:20 CST 2005
#
#**********************************************************************




MACRO INVCKNHD
  PIN I
   AntennaPartialMetalArea                    0.256000 LAYER metal1 ;
   AntennaGateArea                            1.310400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.531140 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    3.341600 LAYER metal1 ;
   AntennaDiffArea                            2.184000 LAYER metal1 ;
  END O

END INVCKNHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:25 CST 2005
#
#**********************************************************************




MACRO INVCKQHD
  PIN I
   AntennaPartialMetalArea                    0.254400 LAYER metal1 ;
   AntennaGateArea                            2.959200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.470941 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   10.476400 LAYER metal1 ;
   AntennaDiffArea                            4.932000 LAYER metal1 ;
  END O

END INVCKQHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:30 CST 2005
#
#**********************************************************************




MACRO INVDHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.883775 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.325200 LAYER metal1 ;
   AntennaDiffArea                            0.516800 LAYER metal1 ;
  END O

END INVDHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:35 CST 2005
#
#**********************************************************************




MACRO INVGHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.284444 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.392400 LAYER metal1 ;
   AntennaDiffArea                            0.720000 LAYER metal1 ;
  END O

END INVGHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:40 CST 2005
#
#**********************************************************************




MACRO INVHHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.451200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.429967 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.968000 LAYER metal1 ;
   AntennaDiffArea                            1.278400 LAYER metal1 ;
  END O

END INVHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:45 CST 2005
#
#**********************************************************************




MACRO INVIHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.561600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.329062 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.731200 LAYER metal1 ;
   AntennaDiffArea                            1.154400 LAYER metal1 ;
  END O

END INVIHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:50 CST 2005
#
#**********************************************************************




MACRO INVJHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.676800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.397161 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.728000 LAYER metal1 ;
   AntennaDiffArea                            1.391200 LAYER metal1 ;
  END O

END INVJHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:16:55 CST 2005
#
#**********************************************************************




MACRO INVKHD
  PIN I
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.902400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.193263 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.724800 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END INVKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:00 CST 2005
#
#**********************************************************************




MACRO INVLHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            1.128000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.141845 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.208000 LAYER metal1 ;
   AntennaDiffArea                            2.143200 LAYER metal1 ;
  END O

END INVLHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:05 CST 2005
#
#**********************************************************************




MACRO INVMHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            1.353600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.101653 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    1.208000 LAYER metal1 ;
   AntennaDiffArea                            2.256000 LAYER metal1 ;
  END O

END INVMHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:10 CST 2005
#
#**********************************************************************




MACRO INVNHD
  PIN I
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            1.804800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.131210 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    2.074800 LAYER metal1 ;
   AntennaDiffArea                            3.008000 LAYER metal1 ;
  END O

END INVNHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:15 CST 2005
#
#**********************************************************************




MACRO INVQHD
  PIN I
   AntennaPartialMetalArea                    0.326000 LAYER metal1 ;
   AntennaGateArea                            4.512000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.242908 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                   11.772000 LAYER metal1 ;
   AntennaDiffArea                            7.520000 LAYER metal1 ;
  END O

END INVQHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:20 CST 2005
#
#**********************************************************************




MACRO INVTCHD
  PIN E
   AntennaPartialMetalArea                    0.342000 LAYER metal1 ;
   AntennaGateArea                            0.152400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.151116 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.122000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.114030 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.395200 LAYER metal1 ;
   AntennaDiffArea                            0.516800 LAYER metal1 ;
  END O

END INVTCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:26 CST 2005
#
#**********************************************************************




MACRO INVTEHD
  PIN E
   AntennaPartialMetalArea                    0.135200 LAYER metal1 ;
   AntennaGateArea                            0.237600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.471376 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.674800 LAYER metal1 ;
   AntennaGateArea                            0.381600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.958846 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.384000 LAYER metal1 ;
   AntennaDiffArea                            0.952000 LAYER metal1 ;
  END O

END INVTEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:32 CST 2005
#
#**********************************************************************




MACRO INVTHHD
  PIN E
   AntennaPartialMetalArea                    0.391200 LAYER metal1 ;
   AntennaGateArea                            0.250800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.502821 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.143600 LAYER metal1 ;
   AntennaGateArea                            0.084000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.714286 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.580000 LAYER metal1 ;
   AntennaDiffArea                            1.008000 LAYER metal1 ;
  END O

END INVTHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:38 CST 2005
#
#**********************************************************************




MACRO INVTKHD
  PIN E
   AntennaPartialMetalArea                    0.416800 LAYER metal1 ;
   AntennaGateArea                            0.273600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.509258 LAYER metal1 ; 
  END E

  PIN I
   AntennaPartialMetalArea                    0.143600 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.065215 LAYER metal1 ; 
  END I

  PIN O
   AntennaPartialMetalArea                    0.808000 LAYER metal1 ;
   AntennaDiffArea                            1.344000 LAYER metal1 ;
  END O

END INVTKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:44 CST 2005
#
#**********************************************************************




MACRO MAO222CHD
  PIN A1
   AntennaPartialMetalArea                    0.140000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.283338 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.816662 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.813600 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.594440 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.319600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END MAO222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:49 CST 2005
#
#**********************************************************************




MACRO MAO222EHD
  PIN A1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.916670 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.377600 LAYER metal1 ;
   AntennaGateArea                            0.384000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.004167 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.687200 LAYER metal1 ;
   AntennaGateArea                            0.355200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.318625 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.319600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END MAO222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:17:55 CST 2005
#
#**********************************************************************




MACRO MAO222HHD
  PIN A1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814810 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.377600 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.892596 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.687200 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.996299 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.364000 LAYER metal1 ;
   AntennaDiffArea                            0.789600 LAYER metal1 ;
  END O

END MAO222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:00 CST 2005
#
#**********************************************************************




MACRO MAO222KHD
  PIN A1
   AntennaPartialMetalArea                    0.140000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.283338 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.816662 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.813600 LAYER metal1 ;
   AntennaGateArea                            0.288000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.594440 LAYER metal1 ; 
  END C1

  PIN O
   AntennaPartialMetalArea                    0.738000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END MAO222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:05 CST 2005
#
#**********************************************************************




MACRO MAOI1CHD
  PIN A1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.007097 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709224 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.738891 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.388890 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.574400 LAYER metal1 ;
   AntennaDiffArea                            0.892800 LAYER metal1 ;
  END O

END MAOI1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:10 CST 2005
#
#**********************************************************************




MACRO MAOI1EHD
  PIN A1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.864583 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.500000 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.523080 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.394872 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.367200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END MAOI1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:16 CST 2005
#
#**********************************************************************




MACRO MAOI1HHD
  PIN A1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.093333 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.860000 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.945098 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.890196 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.565600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END MAOI1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:21 CST 2005
#
#**********************************************************************




MACRO MAOI1KHD
  PIN A1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.007097 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709224 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.738891 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.388890 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.944000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END MAOI1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:26 CST 2005
#
#**********************************************************************




MACRO MOAI1CHD
  PIN A1
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785182 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785190 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.113333 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.880000 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.724800 LAYER metal1 ;
   AntennaDiffArea                            0.730000 LAYER metal1 ;
  END O

END MOAI1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:32 CST 2005
#
#**********************************************************************




MACRO MOAI1EHD
  PIN A1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.661111 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.466670 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008330 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.212500 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.421600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END MOAI1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:37 CST 2005
#
#**********************************************************************




MACRO MOAI1HHD
  PIN A1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.661111 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.466670 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837034 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.940740 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.392400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END MOAI1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:42 CST 2005
#
#**********************************************************************




MACRO MOAI1KHD
  PIN A1
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785182 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785190 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.113333 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.880000 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.736000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END MOAI1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:47 CST 2005
#
#**********************************************************************




MACRO MUX2CHD
  PIN A
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.098400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.772359 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.098400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.065039 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    0.380600 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.962366 LAYER metal1 ; 
  END S

END MUX2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:52 CST 2005
#
#**********************************************************************




MACRO MUX2EHD
  PIN A
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.114000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.403511 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.114000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.529826 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    0.481800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.612289 LAYER metal1 ; 
  END S

END MUX2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:18:57 CST 2005
#
#**********************************************************************




MACRO MUX2HHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792589 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740743 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    0.584000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.651200 LAYER metal1 ;
   AntennaGateArea                            0.242400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.935181 LAYER metal1 ; 
  END S

END MUX2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:02 CST 2005
#
#**********************************************************************




MACRO MUX2KHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.792589 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.740743 LAYER metal1 ; 
  END B

  PIN O
   AntennaPartialMetalArea                    1.000000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.651200 LAYER metal1 ;
   AntennaGateArea                            0.249600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.935186 LAYER metal1 ; 
  END S

END MUX2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:07 CST 2005
#
#**********************************************************************




MACRO MUX3CHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.241023 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.564106 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.160000 LAYER metal1 ;
   AntennaGateArea                            0.098400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.845524 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    0.378400 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.103200 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.043012 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.962364 LAYER metal1 ; 
  END S1

END MUX3CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:11 CST 2005
#
#**********************************************************************




MACRO MUX3EHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.949016 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.031375 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.160000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.133329 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    0.378400 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.103200 LAYER metal1 ;
   AntennaGateArea                            0.153600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.947915 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.516906 LAYER metal1 ; 
  END S1

END MUX3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:17 CST 2005
#
#**********************************************************************




MACRO MUX3HHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758867 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709224 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.025638 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    0.584000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.651200 LAYER metal1 ;
   AntennaGateArea                            0.273600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.935183 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.622400 LAYER metal1 ;
   AntennaGateArea                            0.273600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.935186 LAYER metal1 ; 
  END S1

END MUX3HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:22 CST 2005
#
#**********************************************************************




MACRO MUX3KHD
  PIN A
   AntennaPartialMetalArea                    0.137600 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.922221 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.432000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.805556 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709222 LAYER metal1 ; 
  END C

  PIN O
   AntennaPartialMetalArea                    1.000000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.750400 LAYER metal1 ;
   AntennaGateArea                            0.273600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.935190 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.636800 LAYER metal1 ;
   AntennaGateArea                            0.273600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.935185 LAYER metal1 ; 
  END S1

END MUX3KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:27 CST 2005
#
#**********************************************************************




MACRO MUX4CHD
  PIN A
   AntennaPartialMetalArea                    0.136000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251285 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.205126 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.150001 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.056413 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.309200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.151600 LAYER metal1 ;
   AntennaGateArea                            0.285600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.291318 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.446761 LAYER metal1 ; 
  END S1

END MUX4CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:32 CST 2005
#
#**********************************************************************




MACRO MUX4EHD
  PIN A
   AntennaPartialMetalArea                    0.136000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954167 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.979170 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.150001 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833333 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.309200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.151600 LAYER metal1 ;
   AntennaGateArea                            0.369600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.231597 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.782519 LAYER metal1 ; 
  END S1

END MUX4EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:37 CST 2005
#
#**********************************************************************




MACRO MUX4HHD
  PIN A
   AntennaPartialMetalArea                    0.136000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954167 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.979170 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.150001 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833333 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.309200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.151600 LAYER metal1 ;
   AntennaGateArea                            0.415200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.766855 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.217200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.333336 LAYER metal1 ; 
  END S1

END MUX4HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:42 CST 2005
#
#**********************************************************************




MACRO MUX4KHD
  PIN A
   AntennaPartialMetalArea                    0.136000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090476 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.119046 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.186443 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.952382 LAYER metal1 ; 
  END D

  PIN O
   AntennaPartialMetalArea                    0.944000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.151600 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.601239 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.112400 LAYER metal1 ;
   AntennaGateArea                            0.200400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.421162 LAYER metal1 ; 
  END S1

END MUX4KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:48 CST 2005
#
#**********************************************************************




MACRO MUX5EHD
  PIN A
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.174361 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.140000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.282054 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.150001 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.071793 LAYER metal1 ; 
  END D

  PIN E
   AntennaPartialMetalArea                    0.172400 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.246152 LAYER metal1 ; 
  END E

  PIN O
   AntennaPartialMetalArea                    0.365200 LAYER metal1 ;
   AntennaDiffArea                            0.733200 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.151600 LAYER metal1 ;
   AntennaGateArea                            0.348000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.342528 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.150000 LAYER metal1 ;
   AntennaGateArea                            0.194400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.553495 LAYER metal1 ; 
  END S1

  PIN S2
   AntennaPartialMetalArea                    0.189200 LAYER metal1 ;
   AntennaGateArea                            0.194400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.471189 LAYER metal1 ; 
  END S2

END MUX5EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:53 CST 2005
#
#**********************************************************************




MACRO MUXB2BHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.266662 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.579486 LAYER metal1 ; 
  END B

  PIN EB
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.138000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.463767 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.535200 LAYER metal1 ;
   AntennaDiffArea                            0.412000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.817948 LAYER metal1 ; 
  END S

END MUXB2BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:19:59 CST 2005
#
#**********************************************************************




MACRO MUXB2CHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.983333 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.395239 LAYER metal1 ; 
  END B

  PIN EB
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.933329 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.529200 LAYER metal1 ;
   AntennaDiffArea                            0.520000 LAYER metal1 ;
  END O

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.171600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.582751 LAYER metal1 ; 
  END S

END MUXB2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:04 CST 2005
#
#**********************************************************************




MACRO MUXB4CHD
  PIN A
   AntennaPartialMetalArea                    0.136000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839213 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.921571 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.150001 LAYER metal1 ; 
  END C

  PIN D
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784316 LAYER metal1 ; 
  END D

  PIN EB
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.254025 LAYER metal1 ; 
  END EB

  PIN O
   AntennaPartialMetalArea                    0.463600 LAYER metal1 ;
   AntennaDiffArea                            0.583000 LAYER metal1 ;
  END O

  PIN S0
   AntennaPartialMetalArea                    0.151600 LAYER metal1 ;
   AntennaGateArea                            0.326400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718139 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.852087 LAYER metal1 ; 
  END S1

END MUXB4CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:09 CST 2005
#
#**********************************************************************




MACRO MXL2CHD
  PIN A
   AntennaPartialMetalArea                    0.126400 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784312 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.126400 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839212 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    0.637600 LAYER metal1 ;
   AntennaDiffArea                            0.876000 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.290400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.260333 LAYER metal1 ; 
  END S

END MXL2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:15 CST 2005
#
#**********************************************************************




MACRO MXL2EHD
  PIN A
   AntennaPartialMetalArea                    0.116800 LAYER metal1 ;
   AntennaGateArea                            0.098400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.772358 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.098400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.065039 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    0.457600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.962366 LAYER metal1 ; 
  END S

END MXL2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:20 CST 2005
#
#**********************************************************************




MACRO MXL2HHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.952382 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.395239 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    0.564000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.810258 LAYER metal1 ; 
  END S

END MXL2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:26 CST 2005
#
#**********************************************************************




MACRO MXL2KHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.952382 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.395239 LAYER metal1 ; 
  END B

  PIN OB
   AntennaPartialMetalArea                    0.980000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END OB

  PIN S
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.171600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.582751 LAYER metal1 ; 
  END S

END MXL2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:31 CST 2005
#
#**********************************************************************




MACRO MXL3EHD
  PIN A
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.241023 LAYER metal1 ; 
  END A

  PIN B
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.564106 LAYER metal1 ; 
  END B

  PIN C
   AntennaPartialMetalArea                    0.160000 LAYER metal1 ;
   AntennaGateArea                            0.098400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.845524 LAYER metal1 ; 
  END C

  PIN OB
   AntennaPartialMetalArea                    0.468600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END OB

  PIN S0
   AntennaPartialMetalArea                    0.103200 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.043012 LAYER metal1 ; 
  END S0

  PIN S1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.962364 LAYER metal1 ; 
  END S1

END MXL3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:37 CST 2005
#
#**********************************************************************




MACRO ND2CHD
  PIN I1
   AntennaPartialMetalArea                    0.175600 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.485877 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.310815 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.451200 LAYER metal1 ;
   AntennaDiffArea                            0.437200 LAYER metal1 ;
  END O

END ND2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:42 CST 2005
#
#**********************************************************************




MACRO ND2DHD
  PIN I1
   AntennaPartialMetalArea                    0.175600 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.308460 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.182929 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.451200 LAYER metal1 ;
   AntennaDiffArea                            0.501200 LAYER metal1 ;
  END O

END ND2DHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:47 CST 2005
#
#**********************************************************************




MACRO ND2HHD
  PIN I1
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            0.408000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.852943 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.451200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.771281 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.869600 LAYER metal1 ;
   AntennaDiffArea                            1.116000 LAYER metal1 ;
  END O

END ND2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:52 CST 2005
#
#**********************************************************************




MACRO ND2KHD
  PIN I1
   AntennaPartialMetalArea                    0.818400 LAYER metal1 ;
   AntennaGateArea                            0.777600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.509801 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.799200 LAYER metal1 ;
   AntennaGateArea                            0.806400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.990199 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    2.715200 LAYER metal1 ;
   AntennaDiffArea                            2.342400 LAYER metal1 ;
  END O

END ND2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:20:57 CST 2005
#
#**********************************************************************




MACRO ND3CHD
  PIN I1
   AntennaPartialMetalArea                    0.237600 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.198315 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.856535 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.215200 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.869199 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.838400 LAYER metal1 ;
   AntennaDiffArea                            0.813600 LAYER metal1 ;
  END O

END ND3CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:02 CST 2005
#
#**********************************************************************




MACRO ND3EHD
  PIN I1
   AntennaPartialMetalArea                    0.162000 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.146670 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.151200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.580000 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.722800 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.324442 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.246400 LAYER metal1 ;
   AntennaDiffArea                            1.144000 LAYER metal1 ;
  END O

END ND3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:06 CST 2005
#
#**********************************************************************




MACRO ND3HHD
  PIN I1
   AntennaPartialMetalArea                    0.269600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.290478 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.095235 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.215200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.109528 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.684000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END ND3HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:11 CST 2005
#
#**********************************************************************




MACRO ND4CHD
  PIN I1
   AntennaPartialMetalArea                    0.156000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.988091 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.321430 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.163600 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.345236 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.129600 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.845239 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.348800 LAYER metal1 ;
   AntennaDiffArea                            0.416800 LAYER metal1 ;
  END O

END ND4CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:16 CST 2005
#
#**********************************************************************




MACRO ND4EHD
  PIN I1
   AntennaPartialMetalArea                    0.156000 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.489580 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.906253 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.163600 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.739582 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.129600 LAYER metal1 ;
   AntennaGateArea                            0.076800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.302080 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.558400 LAYER metal1 ;
   AntennaDiffArea                            0.699200 LAYER metal1 ;
  END O

END ND4EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:21 CST 2005
#
#**********************************************************************




MACRO ND4HHD
  PIN I1
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.634925 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.190480 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.163600 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.611114 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.129600 LAYER metal1 ;
   AntennaGateArea                            0.100800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.277776 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.594400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END ND4HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:26 CST 2005
#
#**********************************************************************




MACRO ND4KHD
  PIN I1
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.073333 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.760003 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.163600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.093337 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.129600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.813330 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.544000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END ND4KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:31 CST 2005
#
#**********************************************************************




MACRO ND5EHD
  PIN I1
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.415462 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.122400 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.178740 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.178741 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.181600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.485718 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.188800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.085710 LAYER metal1 ; 
  END I5

  PIN O
   AntennaPartialMetalArea                    0.869600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END ND5EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:36 CST 2005
#
#**********************************************************************




MACRO ND5HHD
  PIN I1
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.536231 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.196800 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.144924 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.180000 LAYER metal1 ;
   AntennaGateArea                            0.165600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.178743 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.181600 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.405407 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.188800 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.027027 LAYER metal1 ; 
  END I5

  PIN O
   AntennaPartialMetalArea                    0.698200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END ND5HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:41 CST 2005
#
#**********************************************************************




MACRO ND6EHD
  PIN I1
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.525250 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.142400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277780 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.120000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.277774 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.172800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.423611 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.249999 LAYER metal1 ; 
  END I5

  PIN I6
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.303026 LAYER metal1 ; 
  END I6

  PIN O
   AntennaPartialMetalArea                    0.553600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END ND6EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:47 CST 2005
#
#**********************************************************************




MACRO ND8DHD
  PIN I1
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.125004 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.206400 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.954545 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.160800 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.212123 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.628784 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.155200 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.946973 LAYER metal1 ; 
  END I5

  PIN I6
   AntennaPartialMetalArea                    0.177600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.636362 LAYER metal1 ; 
  END I6

  PIN I7
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.310604 LAYER metal1 ; 
  END I7

  PIN I8
   AntennaPartialMetalArea                    0.155200 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.685603 LAYER metal1 ; 
  END I8

  PIN O
   AntennaPartialMetalArea                    0.634000 LAYER metal1 ;
   AntennaDiffArea                            0.619200 LAYER metal1 ;
  END O

END ND8DHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:21:53 CST 2005
#
#**********************************************************************




MACRO NR2BHD
  PIN I1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.138000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.918842 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.138000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.428981 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.485600 LAYER metal1 ;
   AntennaDiffArea                            0.412000 LAYER metal1 ;
  END O

END NR2BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:01 CST 2005
#
#**********************************************************************




MACRO NR2CHD
  PIN I1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.031377 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.896935 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.422400 LAYER metal1 ;
   AntennaDiffArea                            0.713200 LAYER metal1 ;
  END O

END NR2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:08 CST 2005
#
#**********************************************************************




MACRO NR2EHD
  PIN I1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.055554 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.606800 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.302224 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.204000 LAYER metal1 ;
   AntennaDiffArea                            1.260000 LAYER metal1 ;
  END O

END NR2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:13 CST 2005
#
#**********************************************************************




MACRO NR2GHD
  PIN I1
   AntennaPartialMetalArea                    0.650000 LAYER metal1 ;
   AntennaGateArea                            0.528000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.166669 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.584800 LAYER metal1 ;
   AntennaGateArea                            0.528000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.473334 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.321600 LAYER metal1 ;
   AntennaDiffArea                            1.481600 LAYER metal1 ;
  END O

END NR2GHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:19 CST 2005
#
#**********************************************************************




MACRO NR2IHD
  PIN I1
   AntennaPartialMetalArea                    1.018400 LAYER metal1 ;
   AntennaGateArea                            0.844800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.273338 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.852400 LAYER metal1 ;
   AntennaGateArea                            0.844800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.300004 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.667200 LAYER metal1 ;
   AntennaDiffArea                            2.146400 LAYER metal1 ;
  END O

END NR2IHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:25 CST 2005
#
#**********************************************************************




MACRO NR3BHD
  PIN I1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.464644 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.464647 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.343434 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.808000 LAYER metal1 ;
   AntennaDiffArea                            0.576800 LAYER metal1 ;
  END O

END NR3BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:31 CST 2005
#
#**********************************************************************




MACRO NR3EHD
  PIN I1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.625646 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.179483 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.241028 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.375200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END NR3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:36 CST 2005
#
#**********************************************************************




MACRO NR3HHD
  PIN I1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.625646 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.179483 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.241028 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.427200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END NR3HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:41 CST 2005
#
#**********************************************************************




MACRO NR4CHD
  PIN I1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.083331 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.287882 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.280301 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.977271 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.333200 LAYER metal1 ;
   AntennaDiffArea                            0.392000 LAYER metal1 ;
  END O

END NR4CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:46 CST 2005
#
#**********************************************************************




MACRO NR4EHD
  PIN I1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.083331 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.287882 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.280301 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.977271 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.395200 LAYER metal1 ;
   AntennaDiffArea                            0.658000 LAYER metal1 ;
  END O

END NR4EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:51 CST 2005
#
#**********************************************************************




MACRO NR4HHD
  PIN I1
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.083331 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.287882 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.280301 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.120800 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.977271 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.462400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END NR4HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:22:57 CST 2005
#
#**********************************************************************




MACRO NR5EHD
  PIN I1
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570617 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.536721 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.858759 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.163200 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.969695 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.969702 LAYER metal1 ; 
  END I5

  PIN O
   AntennaPartialMetalArea                    0.416000 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END NR5EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:02 CST 2005
#
#**********************************************************************




MACRO NR6EHD
  PIN I1
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570622 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.536721 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.858759 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.166400 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.468929 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.116000 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.468931 LAYER metal1 ; 
  END I5

  PIN I6
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.807911 LAYER metal1 ; 
  END I6

  PIN O
   AntennaPartialMetalArea                    0.416000 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END NR6EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:09 CST 2005
#
#**********************************************************************




MACRO NR8EHD
  PIN I1
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.515151 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.045451 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.098489 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.992421 LAYER metal1 ; 
  END I4

  PIN I5
   AntennaPartialMetalArea                    0.126400 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.227270 LAYER metal1 ; 
  END I5

  PIN I6
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.772732 LAYER metal1 ; 
  END I6

  PIN I7
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.954543 LAYER metal1 ; 
  END I7

  PIN I8
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.803032 LAYER metal1 ; 
  END I8

  PIN O
   AntennaPartialMetalArea                    0.656000 LAYER metal1 ;
   AntennaDiffArea                            0.884000 LAYER metal1 ;
  END O

END NR8EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:15 CST 2005
#
#**********************************************************************




MACRO OA112CHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.108000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.103700 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.108000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.137037 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251282 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.502564 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.431600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OA112CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:21 CST 2005
#
#**********************************************************************




MACRO OA112EHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287183 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.310253 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837038 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.018516 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.404800 LAYER metal1 ;
   AntennaDiffArea                            0.614000 LAYER metal1 ;
  END O

END OA112EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:28 CST 2005
#
#**********************************************************************




MACRO OA112HHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.982218 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.002222 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837038 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.018516 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.690400 LAYER metal1 ;
   AntennaDiffArea                            1.309600 LAYER metal1 ;
  END O

END OA112HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:33 CST 2005
#
#**********************************************************************




MACRO OA112KHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.982218 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.002222 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837038 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.018516 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.038400 LAYER metal1 ;
   AntennaDiffArea                            2.091600 LAYER metal1 ;
  END O

END OA112KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:38 CST 2005
#
#**********************************************************************




MACRO OA12CHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.084000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.461903 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.131200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.426667 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.633330 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.394000 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OA12CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:43 CST 2005
#
#**********************************************************************




MACRO OA12EHD
  PIN A1
   AntennaPartialMetalArea                    0.144000 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.884851 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.131200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.447618 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.395240 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.414000 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OA12EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:48 CST 2005
#
#**********************************************************************




MACRO OA12HHD
  PIN A1
   AntennaPartialMetalArea                    0.153200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.247615 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.127200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.909801 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.031369 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.736800 LAYER metal1 ;
   AntennaDiffArea                            1.278400 LAYER metal1 ;
  END O

END OA12HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:54 CST 2005
#
#**********************************************************************




MACRO OA12KHD
  PIN A1
   AntennaPartialMetalArea                    0.153200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.091663 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.127200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.859261 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.974076 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.028800 LAYER metal1 ;
   AntennaDiffArea                            2.030400 LAYER metal1 ;
  END O

END OA12KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:23:59 CST 2005
#
#**********************************************************************




MACRO OA13CHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.566667 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.561107 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.527781 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.566663 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.421200 LAYER metal1 ;
   AntennaDiffArea                            0.398800 LAYER metal1 ;
  END O

END OA13CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:05 CST 2005
#
#**********************************************************************




MACRO OA13EHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.503033 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.920830 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.895833 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.895833 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.421200 LAYER metal1 ;
   AntennaDiffArea                            0.669200 LAYER metal1 ;
  END O

END OA13EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:11 CST 2005
#
#**********************************************************************




MACRO OA13HHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.925928 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837038 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785184 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.468000 LAYER metal1 ;
   AntennaDiffArea                            0.762000 LAYER metal1 ;
  END O

END OA13HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:18 CST 2005
#
#**********************************************************************




MACRO OA13KHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.925928 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837038 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785184 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785190 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.695200 LAYER metal1 ;
   AntennaDiffArea                            1.584000 LAYER metal1 ;
  END O

END OA13KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:24 CST 2005
#
#**********************************************************************




MACRO OA2222CHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.507691 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.210261 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251286 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.502564 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.507695 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.210254 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251278 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.179491 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.689600 LAYER metal1 ;
   AntennaDiffArea                            0.546000 LAYER metal1 ;
  END O

END OA2222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:31 CST 2005
#
#**********************************************************************




MACRO OA2222EHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.035290 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.807840 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839218 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.031369 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.035298 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.807838 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839214 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784310 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.960800 LAYER metal1 ;
   AntennaDiffArea                            1.240000 LAYER metal1 ;
  END O

END OA2222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:37 CST 2005
#
#**********************************************************************




MACRO OA2222HHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.035290 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.807840 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839218 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.031369 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.035298 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.807838 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839214 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784310 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    1.715600 LAYER metal1 ;
   AntennaDiffArea                            2.136000 LAYER metal1 ;
  END O

END OA2222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:44 CST 2005
#
#**********************************************************************




MACRO OA222CHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.261907 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.261907 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.411903 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.261907 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.354763 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.407146 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.431600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OA222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:51 CST 2005
#
#**********************************************************************




MACRO OA222EHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.953701 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837034 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066215 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.949999 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.440400 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OA222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:24:58 CST 2005
#
#**********************************************************************




MACRO OA222HHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.953701 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837034 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066215 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.949999 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.702400 LAYER metal1 ;
   AntennaDiffArea                            1.308400 LAYER metal1 ;
  END O

END OA222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:04 CST 2005
#
#**********************************************************************




MACRO OA222KHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837040 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.953701 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.837034 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066215 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.949999 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.050400 LAYER metal1 ;
   AntennaDiffArea                            2.090400 LAYER metal1 ;
  END O

END OA222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:11 CST 2005
#
#**********************************************************************




MACRO OA22CHD
  PIN A1
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.896970 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.630305 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.678787 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.975761 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.369600 LAYER metal1 ;
   AntennaDiffArea                            0.404800 LAYER metal1 ;
  END O

END OA22CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:17 CST 2005
#
#**********************************************************************




MACRO OA22EHD
  PIN A1
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.124441 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.928888 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.964446 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.182227 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.424800 LAYER metal1 ;
   AntennaDiffArea                            0.631000 LAYER metal1 ;
  END O

END OA22EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:22 CST 2005
#
#**********************************************************************




MACRO OA22HHD
  PIN A1
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.886520 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.730496 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758861 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.715200 LAYER metal1 ;
   AntennaDiffArea                            1.272000 LAYER metal1 ;
  END O

END OA22HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:29 CST 2005
#
#**********************************************************************




MACRO OA22KHD
  PIN A1
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.886520 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.730496 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758861 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.932623 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.016000 LAYER metal1 ;
   AntennaDiffArea                            2.042800 LAYER metal1 ;
  END O

END OA22KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:35 CST 2005
#
#**********************************************************************




MACRO OAI112BHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.327782 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.536108 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954170 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.700000 LAYER metal1 ;
   AntennaDiffArea                            0.856000 LAYER metal1 ;
  END O

END OAI112BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:40 CST 2005
#
#**********************************************************************




MACRO OAI112EHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.108000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.103700 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.108000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.137037 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251282 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.502564 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.334000 LAYER metal1 ;
   AntennaDiffArea                            0.709200 LAYER metal1 ;
  END O

END OAI112EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:47 CST 2005
#
#**********************************************************************




MACRO OAI112HHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.327782 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.352778 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954170 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.460000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OAI112HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:53 CST 2005
#
#**********************************************************************




MACRO OAI112KHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.327782 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.352778 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954170 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.736000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OAI112KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:25:59 CST 2005
#
#**********************************************************************




MACRO OAI12CHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.352778 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954163 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.472800 LAYER metal1 ;
   AntennaDiffArea                            0.604000 LAYER metal1 ;
  END O

END OAI12CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:06 CST 2005
#
#**********************************************************************




MACRO OAI12EHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.838333 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.251286 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.502564 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.308800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OAI12EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:12 CST 2005
#
#**********************************************************************




MACRO OAI12HHD
  PIN A1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.612126 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.208886 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.302227 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.528000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OAI12HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:18 CST 2005
#
#**********************************************************************




MACRO OAI12KHD
  PIN A1
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.144000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.352778 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.954163 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.736000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OAI12KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:25 CST 2005
#
#**********************************************************************




MACRO OAI13BHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.943333 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.048886 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.022226 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.302227 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.513200 LAYER metal1 ;
   AntennaDiffArea                            0.565000 LAYER metal1 ;
  END O

END OAI13BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:31 CST 2005
#
#**********************************************************************




MACRO OAI13EHD
  PIN A1
   AntennaPartialMetalArea                    0.143600 LAYER metal1 ;
   AntennaGateArea                            0.108000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.085180 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.121200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.793938 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.757577 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.139391 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.434000 LAYER metal1 ;
   AntennaDiffArea                            0.709200 LAYER metal1 ;
  END O

END OAI13EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:40 CST 2005
#
#**********************************************************************




MACRO OAI13HHD
  PIN A1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.248719 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.920833 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.895833 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.528000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OAI13HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:48 CST 2005
#
#**********************************************************************




MACRO OAI13KHD
  PIN A1
   AntennaPartialMetalArea                    0.128800 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.248719 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.920833 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.895833 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.158330 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.736000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OAI13KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:26:56 CST 2005
#
#**********************************************************************




MACRO OAI2222CHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.134614 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.762824 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.814101 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.128202 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.134611 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.762822 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.814103 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.124800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.724354 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.381200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OAI2222CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:27:05 CST 2005
#
#**********************************************************************




MACRO OAI2222EHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328573 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052383 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090477 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.323810 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328570 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052386 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090476 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.023813 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.386800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OAI2222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:27:15 CST 2005
#
#**********************************************************************




MACRO OAI2222HHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328573 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052383 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090477 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.323810 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328570 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052386 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090476 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.023813 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.391600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OAI2222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:27:26 CST 2005
#
#**********************************************************************




MACRO OAI2222KHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328573 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052383 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090477 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.323810 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.328570 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.148800 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052386 LAYER metal1 ; 
  END C2

  PIN D1
   AntennaPartialMetalArea                    0.115200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.090476 LAYER metal1 ; 
  END D1

  PIN D2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.023813 LAYER metal1 ; 
  END D2

  PIN O
   AntennaPartialMetalArea                    0.784000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OAI2222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:27:38 CST 2005
#
#**********************************************************************




MACRO OAI222BHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.210000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.761903 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.210000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.767623 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.210000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.841907 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.210000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.855233 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.159600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.962747 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.210000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.977139 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.739600 LAYER metal1 ;
   AntennaDiffArea                            1.100000 LAYER metal1 ;
  END O

END OAI222BHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:27:48 CST 2005
#
#**********************************************************************




MACRO OAI222EHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.760607 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.760607 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.951515 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.760601 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.878786 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.945450 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.303200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OAI222EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:27:55 CST 2005
#
#**********************************************************************




MACRO OAI222HHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066664 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066664 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.211492 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.066671 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.156324 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.174000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.206899 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.368000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OAI222HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:03 CST 2005
#
#**********************************************************************




MACRO OAI222KHD
  PIN A1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.186000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.965594 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.186000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.965594 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.186000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.101079 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.156800 LAYER metal1 ;
   AntennaGateArea                            0.186000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.965589 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.137200 LAYER metal1 ;
   AntennaGateArea                            0.186000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.049466 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.186000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.096773 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.736000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OAI222KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:12 CST 2005
#
#**********************************************************************




MACRO OAI22CHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.035290 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.807840 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.839218 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.031369 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.422000 LAYER metal1 ;
   AntennaDiffArea                            0.680000 LAYER metal1 ;
  END O

END OAI22CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:22 CST 2005
#
#**********************************************************************




MACRO OAI22EHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287181 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.133332 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.317946 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.425644 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.308800 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OAI22EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:31 CST 2005
#
#**********************************************************************




MACRO OAI22HHD
  PIN A1
   AntennaPartialMetalArea                    0.112000 LAYER metal1 ;
   AntennaGateArea                            0.162000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.276542 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.162000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.128390 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.162000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.306176 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.162000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.409874 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.368000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OAI22HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:39 CST 2005
#
#**********************************************************************




MACRO OAI22KHD
  PIN A1
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.195233 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.134400 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052380 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.123200 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.223807 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.117600 LAYER metal1 ;
   AntennaGateArea                            0.168000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.323810 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.736000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OAI22KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:48 CST 2005
#
#**********************************************************************




MACRO OR2B1CHD
  PIN B1
   AntennaPartialMetalArea                    0.113200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.482049 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.855556 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.473600 LAYER metal1 ;
   AntennaDiffArea                            0.548000 LAYER metal1 ;
  END O

END OR2B1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:28:54 CST 2005
#
#**********************************************************************




MACRO OR2B1EHD
  PIN B1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.722226 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.113200 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.813337 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.365200 LAYER metal1 ;
   AntennaDiffArea                            0.718400 LAYER metal1 ;
  END O

END OR2B1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:00 CST 2005
#
#**********************************************************************




MACRO OR2B1HHD
  PIN B1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.572226 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.113200 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.358451 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.573000 LAYER metal1 ;
   AntennaDiffArea                            0.864800 LAYER metal1 ;
  END O

END OR2B1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:07 CST 2005
#
#**********************************************************************




MACRO OR2B1KHD
  PIN B1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.108000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.692594 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.118800 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.194440 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.981400 LAYER metal1 ;
   AntennaDiffArea                            1.512800 LAYER metal1 ;
  END O

END OR2B1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:14 CST 2005
#
#**********************************************************************




MACRO OR2CHD
  PIN I1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.280303 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.481062 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.381200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OR2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:22 CST 2005
#
#**********************************************************************




MACRO OR2EHD
  PIN I1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.653333 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.120000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.013333 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.381200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OR2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:29 CST 2005
#
#**********************************************************************




MACRO OR2HHD
  PIN I1
   AntennaPartialMetalArea                    0.112800 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.260274 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.703198 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.448400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OR2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:36 CST 2005
#
#**********************************************************************




MACRO OR2KHD
  PIN I1
   AntennaPartialMetalArea                    0.561600 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.393520 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.247684 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.080000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END OR2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:44 CST 2005
#
#**********************************************************************




MACRO OR3B1CHD
  PIN B1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.688886 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.299439 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.135600 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.299433 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.375200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OR3B1CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:51 CST 2005
#
#**********************************************************************




MACRO OR3B1EHD
  PIN B1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.655556 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.179489 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.135600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.179489 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.375200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OR3B1EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:29:58 CST 2005
#
#**********************************************************************




MACRO OR3B1HHD
  PIN B1
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.255556 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.612000 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.933332 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.461200 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.292305 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.456000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OR3B1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:06 CST 2005
#
#**********************************************************************




MACRO OR3B2CHD
  PIN B1
   AntennaPartialMetalArea                    0.143200 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.930738 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.930736 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.086400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.935185 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.674000 LAYER metal1 ;
   AntennaDiffArea                            0.787600 LAYER metal1 ;
  END O

END OR3B2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:14 CST 2005
#
#**********************************************************************




MACRO OR3B2EHD
  PIN B1
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.088887 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.072000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.788886 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.111200 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.179489 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.375200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OR3B2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:22 CST 2005
#
#**********************************************************************




MACRO OR3B2HHD
  PIN B1
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.484845 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.866668 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.612800 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008337 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.468800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OR3B2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:29 CST 2005
#
#**********************************************************************




MACRO OR3B2KHD
  PIN B1
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.506065 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.107600 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.866668 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.613600 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.015623 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.934400 LAYER metal1 ;
   AntennaDiffArea                            1.524000 LAYER metal1 ;
  END O

END OR3B2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:38 CST 2005
#
#**********************************************************************




MACRO OR3CHD
  PIN I1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.519778 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.757067 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.858758 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.367200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END O

END OR3CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:45 CST 2005
#
#**********************************************************************




MACRO OR3EHD
  PIN I1
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.287182 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.487176 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.156000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.610255 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.367200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END OR3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:52 CST 2005
#
#**********************************************************************




MACRO OR3HHD
  PIN I1
   AntennaPartialMetalArea                    0.645600 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.213329 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.396800 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.333335 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.312000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.928206 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.434400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END O

END OR3HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:30:59 CST 2005
#
#**********************************************************************




MACRO QDBAHEHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.139200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.347696 LAYER metal1 ; 
  END D

  PIN GB
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END GB

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

END QDBAHEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:07 CST 2005
#
#**********************************************************************




MACRO QDBAHHHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783690 LAYER metal1 ; 
  END D

  PIN GB
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.603770 LAYER metal1 ; 
  END GB

  PIN Q
   AntennaPartialMetalArea                    0.326800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

END QDBAHHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:15 CST 2005
#
#**********************************************************************




MACRO QDFFCHD
  PIN CK
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.097777 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.359200 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END Q

END QDFFCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:24 CST 2005
#
#**********************************************************************




MACRO QDFFEHD
  PIN CK
   AntennaPartialMetalArea                    0.144400 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570918 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.419200 LAYER metal1 ;
   AntennaDiffArea                            0.457200 LAYER metal1 ;
  END Q

END QDFFEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:31 CST 2005
#
#**********************************************************************




MACRO QDFFHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570922 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.421600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

END QDFFHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:40 CST 2005
#
#**********************************************************************




MACRO QDFFKHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.808000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

END QDFFKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:47 CST 2005
#
#**********************************************************************




MACRO QDFFRBCHD
  PIN CK
   AntennaPartialMetalArea                    0.149200 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.177782 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.335200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.165600 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.749512 LAYER metal1 ; 
  END RB

END QDFFRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:31:53 CST 2005
#
#**********************************************************************




MACRO QDFFRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.149200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609925 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.243200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.165600 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.702172 LAYER metal1 ; 
  END RB

END QDFFRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:00 CST 2005
#
#**********************************************************************




MACRO QDFFRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.154800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609930 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.310400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

END QDFFRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:07 CST 2005
#
#**********************************************************************




MACRO QDFFRBKHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709217 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.766670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.130400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

END QDFFRBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:15 CST 2005
#
#**********************************************************************




MACRO QDFFRSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634752 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.112497 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.251200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.165000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.317209 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.116400 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.689266 LAYER metal1 ; 
  END SB

END QDFFRSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:22 CST 2005
#
#**********************************************************************




MACRO QDFFRSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634752 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.112497 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.428400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.612744 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.174861 LAYER metal1 ; 
  END SB

END QDFFRSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:30 CST 2005
#
#**********************************************************************




MACRO QDFFSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609932 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.283200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN SB
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.571758 LAYER metal1 ; 
  END SB

END QDFFSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:37 CST 2005
#
#**********************************************************************




MACRO QDFFSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609932 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.141600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.791670 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.415200 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN SB
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.247965 LAYER metal1 ; 
  END SB

END QDFFSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:45 CST 2005
#
#**********************************************************************




MACRO QDFZCHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.128890 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.359200 LAYER metal1 ;
   AntennaDiffArea                            0.358400 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END QDFZCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:32:52 CST 2005
#
#**********************************************************************




MACRO QDFZEHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.429200 LAYER metal1 ;
   AntennaDiffArea                            0.457200 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END QDFZEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:33:14 CST 2005
#
#**********************************************************************




MACRO QDFZHHD
  PIN CK
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.570919 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.393600 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.291669 LAYER metal1 ; 
  END TD

END QDFZHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:33:36 CST 2005
#
#**********************************************************************




MACRO QDFZKHD
  PIN CK
   AntennaPartialMetalArea                    0.119200 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709221 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.808000 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.528989 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.106000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.898809 LAYER metal1 ; 
  END TD

END QDFZKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:33:43 CST 2005
#
#**********************************************************************




MACRO QDFZRBCHD
  PIN CK
   AntennaPartialMetalArea                    0.108000 LAYER metal1 ;
   AntennaGateArea                            0.090000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.311110 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.433200 LAYER metal1 ;
   AntennaDiffArea                            0.401200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.976332 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.746379 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END QDFZRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:33:50 CST 2005
#
#**********************************************************************




MACRO QDFZRBEHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843967 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.310400 LAYER metal1 ;
   AntennaDiffArea                            0.454400 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.202800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.702172 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END QDFZRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:34:13 CST 2005
#
#**********************************************************************




MACRO QDFZRBHHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.843967 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.310400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END QDFZRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:34:34 CST 2005
#
#**********************************************************************




MACRO QDFZRBKHD
  PIN CK
   AntennaPartialMetalArea                    0.124800 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.709219 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.134800 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854705 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    1.130400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.132000 LAYER metal1 ;
   AntennaGateArea                            0.292800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.490440 LAYER metal1 ; 
  END RB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.583329 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.164800 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.023809 LAYER metal1 ; 
  END TD

END QDFZRBKHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:34:42 CST 2005
#
#**********************************************************************




MACRO QDFZRSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.110800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634750 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.918799 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.321600 LAYER metal1 ;
   AntennaDiffArea                            0.555200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.160000 LAYER metal1 ;
   AntennaGateArea                            0.148800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.413981 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.113600 LAYER metal1 ;
   AntennaGateArea                            0.141600 LAYER metal1 ;
   AntennaMaxAreaCAR                          6.689270 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.507249 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.309521 LAYER metal1 ; 
  END TD

END QDFZRSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:34:50 CST 2005
#
#**********************************************************************




MACRO QDFZRSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.110800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.634750 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.918799 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.464000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.108400 LAYER metal1 ;
   AntennaGateArea                            0.244800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.681370 LAYER metal1 ; 
  END RB

  PIN SB
   AntennaPartialMetalArea                    0.133200 LAYER metal1 ;
   AntennaGateArea                            0.146400 LAYER metal1 ;
   AntennaMaxAreaCAR                          7.163934 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.507249 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.309521 LAYER metal1 ; 
  END TD

END QDFZRSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:34:58 CST 2005
#
#**********************************************************************




MACRO QDFZSBEHD
  PIN CK
   AntennaPartialMetalArea                    0.116400 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.609925 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854699 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.243200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN SB
   AntennaPartialMetalArea                    0.104000 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.537038 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.670289 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.404761 LAYER metal1 ; 
  END TD

END QDFZSBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:06 CST 2005
#
#**********************************************************************




MACRO QDFZSBHHD
  PIN CK
   AntennaPartialMetalArea                    0.152800 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.734040 LAYER metal1 ; 
  END CK

  PIN D
   AntennaPartialMetalArea                    0.129200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.854699 LAYER metal1 ; 
  END D

  PIN Q
   AntennaPartialMetalArea                    0.342400 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN SB
   AntennaPartialMetalArea                    0.109600 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.121949 LAYER metal1 ; 
  END SB

  PIN SEL
   AntennaPartialMetalArea                    0.188400 LAYER metal1 ;
   AntennaGateArea                            0.220800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.670289 LAYER metal1 ; 
  END SEL

  PIN TD
   AntennaPartialMetalArea                    0.114000 LAYER metal1 ;
   AntennaGateArea                            0.067200 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.404761 LAYER metal1 ; 
  END TD

END QDFZSBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:14 CST 2005
#
#**********************************************************************




MACRO QDLAHCHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.110400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.688402 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END Q

END QDLAHCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:22 CST 2005
#
#**********************************************************************




MACRO QDLAHEHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.139200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.347696 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

END QDLAHEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:29 CST 2005
#
#**********************************************************************




MACRO QDLAHHHD
  PIN D
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.225600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.783690 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.603770 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.326800 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

END QDLAHHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:36 CST 2005
#
#**********************************************************************




MACRO QDLAHRBCHD
  PIN D
   AntennaPartialMetalArea                    0.163200 LAYER metal1 ;
   AntennaGateArea                            0.177600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.076581 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.091200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.710530 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.380800 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.135200 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976195 LAYER metal1 ; 
  END RB

END QDLAHRBCHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:43 CST 2005
#
#**********************************************************************




MACRO QDLAHRBEHD
  PIN D
   AntennaPartialMetalArea                    0.163200 LAYER metal1 ;
   AntennaGateArea                            0.189600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.008441 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.259600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.135200 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.976195 LAYER metal1 ; 
  END RB

END QDLAHRBEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:51 CST 2005
#
#**********************************************************************




MACRO QDLAHRBHHD
  PIN D
   AntennaPartialMetalArea                    0.205600 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.912699 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.603770 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.368000 LAYER metal1 ;
   AntennaDiffArea                            0.752000 LAYER metal1 ;
  END Q

  PIN RB
   AntennaPartialMetalArea                    0.130000 LAYER metal1 ;
   AntennaGateArea                            0.201600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.063489 LAYER metal1 ; 
  END RB

END QDLAHRBHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:35:58 CST 2005
#
#**********************************************************************




MACRO QDLAHSEHD
  PIN D
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.160800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.054730 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.549997 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.343600 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END Q

  PIN S
   AntennaPartialMetalArea                    0.152000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.348484 LAYER metal1 ; 
  END S

END QDLAHSEHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:05 CST 2005
#
#**********************************************************************




MACRO QDLAHSHHD
  PIN D
   AntennaPartialMetalArea                    0.114800 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.967588 LAYER metal1 ; 
  END D

  PIN G
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.127200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.679250 LAYER metal1 ; 
  END G

  PIN Q
   AntennaPartialMetalArea                    0.643200 LAYER metal1 ;
   AntennaDiffArea                            1.278400 LAYER metal1 ;
  END Q

  PIN S
   AntennaPartialMetalArea                    0.152000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.348484 LAYER metal1 ; 
  END S

END QDLAHSHHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:12 CST 2005
#
#**********************************************************************




MACRO TIE0DHD
  PIN O
   AntennaPartialMetalArea                    0.352400 LAYER metal1 ;
   AntennaDiffArea                            0.238000 LAYER metal1 ;
  END O

END TIE0DHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:18 CST 2005
#
#**********************************************************************




MACRO TIE0HHD
  PIN O
   AntennaPartialMetalArea                    0.428000 LAYER metal1 ;
   AntennaDiffArea                            0.323200 LAYER metal1 ;
  END O

END TIE0HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:25 CST 2005
#
#**********************************************************************




MACRO TIE0KHD
  PIN O
   AntennaPartialMetalArea                    0.824000 LAYER metal1 ;
   AntennaDiffArea                            0.675200 LAYER metal1 ;
  END O

END TIE0KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:32 CST 2005
#
#**********************************************************************




MACRO TIE1DHD
  PIN O
   AntennaPartialMetalArea                    0.351200 LAYER metal1 ;
   AntennaDiffArea                            0.278800 LAYER metal1 ;
  END O

END TIE1DHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:38 CST 2005
#
#**********************************************************************




MACRO TIE1HHD
  PIN O
   AntennaPartialMetalArea                    0.468000 LAYER metal1 ;
   AntennaDiffArea                            0.371200 LAYER metal1 ;
  END O

END TIE1HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:45 CST 2005
#
#**********************************************************************




MACRO TIE1KHD
  PIN O
   AntennaPartialMetalArea                    0.852000 LAYER metal1 ;
   AntennaDiffArea                            0.771200 LAYER metal1 ;
  END O

END TIE1KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:52 CST 2005
#
#**********************************************************************




MACRO XNR2CHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.088800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.621626 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.175200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.817356 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.459200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END XNR2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:36:58 CST 2005
#
#**********************************************************************




MACRO XNR2EHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.088800 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.675676 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.182400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.692986 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.471200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END XNR2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:06 CST 2005
#
#**********************************************************************




MACRO XNR2HHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.117600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.857138 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.230400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.923614 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.536000 LAYER metal1 ;
   AntennaDiffArea                            0.864800 LAYER metal1 ;
  END O

END XNR2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:13 CST 2005
#
#**********************************************************************




MACRO XNR2KHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.999995 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.483200 LAYER metal1 ;
   AntennaGateArea                            0.367200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.362746 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.190400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END XNR2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:20 CST 2005
#
#**********************************************************************




MACRO XNR3CHD
  PIN I1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.112800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.780138 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.278400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.143680 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.184800 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.021643 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.396600 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END XNR3CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:27 CST 2005
#
#**********************************************************************




MACRO XNR3EHD
  PIN I1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.132000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.466663 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.333600 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.328539 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.232800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.017182 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.345400 LAYER metal1 ;
   AntennaDiffArea                            0.714400 LAYER metal1 ;
  END O

END XNR3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:34 CST 2005
#
#**********************************************************************




MACRO XNR4EHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.103200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.162796 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.192000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.408333 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.400003 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.196800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.300813 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.440000 LAYER metal1 ;
   AntennaDiffArea                            0.733200 LAYER metal1 ;
  END O

END XNR4EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:41 CST 2005
#
#**********************************************************************




MACRO XOR2CHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.084000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.771424 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.756800 LAYER metal1 ;
   AntennaGateArea                            0.170400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.047615 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.459200 LAYER metal1 ;
   AntennaDiffArea                            0.384200 LAYER metal1 ;
  END O

END XOR2CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:37:48 CST 2005
#
#**********************************************************************




MACRO XOR2EHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.103200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.162796 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.721600 LAYER metal1 ;
   AntennaGateArea                            0.170400 LAYER metal1 ;
   AntennaMaxAreaCAR                          5.047618 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.471200 LAYER metal1 ;
   AntennaDiffArea                            0.639200 LAYER metal1 ;
  END O

END XOR2EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:38:15 CST 2005
#
#**********************************************************************




MACRO XOR2HHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.199200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.000000 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.734400 LAYER metal1 ;
   AntennaGateArea                            0.237600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.444441 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.536000 LAYER metal1 ;
   AntennaDiffArea                            0.864800 LAYER metal1 ;
  END O

END XOR2HHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:38:36 CST 2005
#
#**********************************************************************




MACRO XOR2KHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.216000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.888894 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.791200 LAYER metal1 ;
   AntennaGateArea                            0.235200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.425924 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.190400 LAYER metal1 ;
   AntennaDiffArea                            1.504000 LAYER metal1 ;
  END O

END XOR2KHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:38:43 CST 2005
#
#**********************************************************************




MACRO XOR3CHD
  PIN I1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.105600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.924239 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.161600 LAYER metal1 ;
   AntennaGateArea                            0.261600 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.400613 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.172800 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.842594 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.387200 LAYER metal1 ;
   AntennaDiffArea                            0.425600 LAYER metal1 ;
  END O

END XOR3CHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:38:50 CST 2005
#
#**********************************************************************




MACRO XOR3EHD
  PIN I1
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.129600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.493826 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.145600 LAYER metal1 ;
   AntennaGateArea                            0.319200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.493730 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.139200 LAYER metal1 ;
   AntennaGateArea                            0.204000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.137257 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.501600 LAYER metal1 ;
   AntennaDiffArea                            0.714400 LAYER metal1 ;
  END O

END XOR3EHD


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Mon May 23 21:38:58 CST 2005
#
#**********************************************************************




MACRO XOR4EHD
  PIN I1
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.400003 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.608889 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.150400 LAYER metal1 ;
   AntennaGateArea                            0.096000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.400003 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.128000 LAYER metal1 ;
   AntennaGateArea                            0.180000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.595559 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.370000 LAYER metal1 ;
   AntennaDiffArea                            0.733200 LAYER metal1 ;
  END O

END XOR4EHD

END LIBRARY
