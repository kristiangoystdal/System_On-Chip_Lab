##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Wed Jan 15 20:07:57 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERcore
  CLASS BLOCK ;
  SIZE 864.000000 BY 363.200000 ;
  FOREIGN BATCHARGERcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN iforcedbat
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.100000 362.680000 0.300000 363.200000 ;
    END
  END iforcedbat
  PIN vsensbat
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 863.700000 362.680000 863.900000 363.200000 ;
    END
  END vsensbat
  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 0.100000 0.000000 0.300000 0.520000 ;
    END
  END vin
  PIN vbattemp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 0.100000 864.000000 0.300000 ;
    END
  END vbattemp
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 362.900000 864.000000 363.100000 ;
    END
  END en
  PIN sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 345.700000 0.000000 345.900000 0.520000 ;
    END
  END sel[3]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 518.500000 0.000000 518.700000 0.520000 ;
    END
  END sel[2]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 691.300000 0.000000 691.500000 0.520000 ;
    END
  END sel[1]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 863.700000 0.000000 863.900000 0.520000 ;
    END
  END sel[0]
  PIN pgnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 172.900000 0.000000 173.100000 0.520000 ;
    END
  END pgnd
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 242.100000 864.000000 242.300000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 121.300000 864.000000 121.500000 ;
    END
  END dgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal2 ;
      RECT 0.500000 362.480000 863.500000 363.200000 ;
      RECT 0.000000 0.720000 864.000000 362.480000 ;
      RECT 691.700000 0.000000 863.500000 0.720000 ;
      RECT 518.900000 0.000000 691.100000 0.720000 ;
      RECT 346.100000 0.000000 518.300000 0.720000 ;
      RECT 173.300000 0.000000 345.500000 0.720000 ;
      RECT 0.500000 0.000000 172.700000 0.720000 ;
    LAYER metal3 ;
      RECT 0.000000 362.700000 863.280000 363.200000 ;
      RECT 0.000000 242.500000 864.000000 362.700000 ;
      RECT 0.000000 241.900000 863.280000 242.500000 ;
      RECT 0.000000 121.700000 864.000000 241.900000 ;
      RECT 0.000000 121.100000 863.280000 121.700000 ;
      RECT 0.000000 0.500000 864.000000 121.100000 ;
      RECT 0.000000 0.000000 863.280000 0.500000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
  END
END BATCHARGERcore

END LIBRARY
