`timescale 1 ns / 10 ps

module BATCHARGERlipo (
    output [63:0] vbat,  // battery voltage (V)
    input [63:0] ibat,  // battery current (A)
    output     [63:0] vtbat     // Voltage proportional to battery temperature: -40ªC to 125ºC are converted in 0V to vref
);

  //-- Default parameters ----------------------------------------------------
  parameter ESR = 0.290;  // Equivalent series resistance (Ohm)
  parameter C = 0.42;  // Capacity (Ah)
  parameter SOC_0 = -0.022;  // Initial state-of-change (0 < SOC < 1))
  // Negative (down to -0.075) can be used for very deeply discharged batteries
  parameter STEP = 10;  // Integration step(ns)
  parameter TIME_STRETCH = 1000000;  // Integration step(ns)

  // Source for LiPo model:
  // Barai, Anup & Widanage, W.D. & Marco, James & Mcgordon, Andrew & Jennings, Paul. (2015). 
  // A study of the open circuit voltage characterization technique and hysteresis assessment of lithium-ion cells. 
  // Journal of Power Sources. 295. 99-107.10.1016/j.jpowsour.2015.06.140.

  parameter a1 = -0.3973;
  parameter b1 = -19.09;
  parameter a2 = 3.549;
  parameter b2 = -0.02769;
  parameter c = 0.7638;
  parameter e = 2.71828;
  parameter rl_ta = 20.0;  // Ambient temperature
  parameter rl_vref = 0.5;  // reference voltage for temperature measurement


  // Thermal heating of battery takes into account 2 contribution: self-heating due to ESR and dissipation due to convection
  //
  //              E_ESR   E_conv
  // T_bat = TA + ----- - ------ , where E_ESR is the integral of the power of heating generated by the ESR 
  //              m * c   m * c 
  //
  //       where E_ESR is the integral of the power of heating generated by the ESR
  //             m: battery mass, for a typical 60 mAh battery m = 2 g
  //             c: thermal capacity of battery (typ. 0.4 J/(gK))
  //
  // E_conv = integral_over_time( h*A*(T_bat - T_A) ),
  //       where h: heat tranfer coefficient of medium around battery (25 W/(m^2 K) for air)
  //             A: contact area (total area of the battery exposed to the air): for a 26x9x3.5mm battery -> A = 0.0007 m^2

  parameter m_bat = 8.8;  // Battery mass in g   
  parameter c_bat = 0.4;  // Battery thermal capacity in J/(gK)
  parameter h = 6;  // Heat tranfer coefficient of medium around battery in W/(m^2 K)
  parameter A = 0.0021;  // Contact area

  //-- Internal signals ------------------------------------------------------
  real rl_vbat;
  real soc;
  real dQ;
  real Q;
  real rl_ibat;
  real rl_ibatdef;  // equal to rl_ibat except if ibat is not defined (in that case rl_ibatdef=0 )    
  real voc;
  real rl_tbat;
  real rl_vtbat;
  real dE_ESR;
  real dE_conv;

  real voc_n;
  real voc_n1;
  real voc_n2;
  real voc_n3;


  // this temperature monitor process is a simplification
  // Real battery temperture is measured using a NTC that requires a series resistor for linearization and a buffer for voltage driving
  initial
    assign rl_vtbat = rl_tbat * rl_vref / 165.0 + 40.0 * rl_vref / 165.0; // converts temperature to voltage: -40 to 125 fitted in the range 0V to vref


  //-- Initial status definition ----------------------------------------------
  initial begin
    soc = SOC_0;
    Q = (C * 60 * 60) * SOC_0;
    voc = a1 * (e ** (b1 * soc)) + a2 * (e ** (b2 * soc)) + c * (soc ** 2);
    voc_n = voc;
    voc_n1 = voc;
    voc_n2 = voc;
    voc_n3 = voc;
    rl_vbat = voc;

    #(STEP / 2);
    rl_tbat = rl_ta;
  end


  //-- Functional --------------------------------------------------------------
  always begin
    #STEP;

    if (^ibat !== 1'bX) rl_ibatdef = rl_ibat;
    else rl_ibatdef = 0;

    dQ = rl_ibat * ((STEP * 1e-9) * TIME_STRETCH);
    Q = Q + dQ;
    soc = Q / (C * 60 * 60);
    voc = a1 * (e ** (b1 * soc)) + a2 * (e ** (b2 * soc)) + c * (soc ** 2);

    rl_vbat = voc;

    // Some settling time
    voc = (voc + voc_n + voc_n1) / 3;
    voc_n = voc;
    voc_n1 = voc_n;

    dE_ESR = (rl_ibat ** 2) * ESR * ((STEP * 1e-9) * TIME_STRETCH);
    dE_conv = h * A * (rl_tbat - rl_ta) * ((STEP * 1e-9) * TIME_STRETCH);
    rl_tbat = rl_tbat + (dE_ESR - dE_conv) / (m_bat * c_bat);
    // rl_tbat = rl_ta;
  end


  //-- Signals conversion ---------------------------------------------------
  initial assign rl_ibat = $bitstoreal(ibat);

  assign vtbat = $realtobits(rl_vtbat);
  assign vbat  = $realtobits(rl_vbat);

endmodule
