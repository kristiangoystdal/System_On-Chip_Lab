##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Thu Jan 16 19:27:24 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BATCHARGERcore
  CLASS BLOCK ;
  SIZE 864.000000 BY 363.200000 ;
  FOREIGN BATCHARGERcore 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN iforcedbat
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 258.900000 864.000000 259.100000 ;
    END
  END iforcedbat
  PIN vsensbat
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 362.900000 864.000000 363.100000 ;
    END
  END vsensbat
  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 699.700000 0.000000 699.900000 0.520000 ;
    END
  END vin
  PIN vbattemp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 154.900000 864.000000 155.100000 ;
    END
  END vbattemp
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 863.480000 50.500000 864.000000 50.700000 ;
    END
  END en
  PIN sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 574.900000 0.000000 575.100000 0.520000 ;
    END
  END sel[3]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 450.100000 0.000000 450.300000 0.520000 ;
    END
  END sel[2]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 325.300000 0.000000 325.500000 0.520000 ;
    END
  END sel[1]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 200.100000 0.000000 200.300000 0.520000 ;
    END
  END sel[0]
  PIN dvdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 399.200000 362.680000 401.200000 363.200000 ;
    END
  END dvdd
  PIN dgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 498.800000 362.680000 500.800000 363.200000 ;
    END
  END dgnd
  PIN pgnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 599.200000 362.680000 601.200000 363.200000 ;
    END
  END pgnd
  OBS
    LAYER metal1 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal2 ;
      RECT 0.000000 0.720000 864.000000 363.200000 ;
      RECT 700.100000 0.000000 864.000000 0.720000 ;
      RECT 575.300000 0.000000 699.500000 0.720000 ;
      RECT 450.500000 0.000000 574.700000 0.720000 ;
      RECT 325.700000 0.000000 449.900000 0.720000 ;
      RECT 200.500000 0.000000 325.100000 0.720000 ;
      RECT 0.000000 0.000000 199.900000 0.720000 ;
    LAYER metal3 ;
      RECT 601.400000 362.700000 863.280000 363.200000 ;
      RECT 601.400000 362.480000 864.000000 362.700000 ;
      RECT 501.000000 362.480000 599.000000 363.200000 ;
      RECT 401.400000 362.480000 498.600000 363.200000 ;
      RECT 0.000000 362.480000 399.000000 363.200000 ;
      RECT 0.000000 259.300000 864.000000 362.480000 ;
      RECT 0.000000 258.700000 863.280000 259.300000 ;
      RECT 0.000000 155.300000 864.000000 258.700000 ;
      RECT 0.000000 154.700000 863.280000 155.300000 ;
      RECT 0.000000 50.900000 864.000000 154.700000 ;
      RECT 0.000000 50.300000 863.280000 50.900000 ;
      RECT 0.000000 0.000000 864.000000 50.300000 ;
    LAYER metal4 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal5 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal6 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal7 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
    LAYER metal8 ;
      RECT 0.000000 0.000000 864.000000 363.200000 ;
  END
END BATCHARGERcore

END LIBRARY
