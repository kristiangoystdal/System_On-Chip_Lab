##
## LEF for PtnCells ;
## created by Innovus v20.11-s130_1 on Sun Dec 19 10:57:57 2021
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO vcobasic
  CLASS BLOCK ;
  SIZE 34.000000 BY 31.200000 ;
  FOREIGN vco 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 9.720000 0.640000 9.880000 ;
    END
  END clk
  PIN vctrl
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 19.320000 0.640000 19.480000 ;
    END
  END vctrl
  PIN avdd
    DIRECTION INOUT ;
#    USE POWER ;
    PORT
      LAYER metal3 ;
        RECT 32.400000 16.000000 34.000000 18.000000 ;
    END
  END avdd
  PIN agnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal3 ;
        RECT 32.400000 4.000000 34.000000 6.000000 ;
    END
  END agnd
 OBS
    LAYER metal1 ;
      RECT 0.000000 21.240000 34.000000 31.200000 ;
      RECT 0.830000 20.760000 34.000000 21.240000 ;
      RECT 0.000000 19.640000 34.000000 20.760000 ;
      RECT 0.830000 19.160000 34.000000 19.640000 ;
      RECT 0.000000 18.040000 34.000000 19.160000 ;
      RECT 0.830000 17.560000 34.000000 18.040000 ;
      RECT 0.000000 16.440000 34.000000 17.560000 ;
      RECT 0.830000 15.960000 34.000000 16.440000 ;
      RECT 0.000000 14.840000 34.000000 15.960000 ;
      RECT 0.830000 14.360000 34.000000 14.840000 ;
      RECT 0.000000 13.240000 34.000000 14.360000 ;
      RECT 0.830000 12.760000 34.000000 13.240000 ;
      RECT 0.000000 11.640000 34.000000 12.760000 ;
      RECT 0.830000 11.160000 34.000000 11.640000 ;
      RECT 0.000000 10.040000 34.000000 11.160000 ;
      RECT 0.830000 9.560000 34.000000 10.040000 ;
      RECT 0.000000 0.000000 34.000000 9.560000 ;
    LAYER metal2 ;
      RECT 0.000000 0.000000 34.000000 31.200000 ;
    LAYER metal3 ;
     RECT 0.000000 18.280000 34.000000 31.200000 ;
     RECT 0.000000 15.720000 32.120000 18.280000 ;
     RECT 0.000000 6.280000 34.000000 15.720000 ;
     RECT 0.000000 3.720000 32.120000 6.280000 ;
     RECT 0.000000 0.000000 34.000000 3.720000 ;
   LAYER metal4 ;
     RECT 0.000000 0.000000 34.000000 31.200000 ;
   LAYER metal5 ;
     RECT 0.000000 0.000000 34.000000 31.200000 ;
   LAYER metal6 ;
     RECT 0.000000 0.000000 34.000000 31.200000 ;
   LAYER metal7 ;
     RECT 0.000000 0.000000 34.000000 31.200000 ;
   LAYER metal8 ;
     RECT 0.000000 0.000000 34.000000 31.200000 ;
 END

END vcobasic

END LIBRARY
