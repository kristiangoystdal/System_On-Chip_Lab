NAMESCASESENSITIVE ON ;
MACRO AN2B1CHD
    CLASS CORE ;
    FOREIGN AN2B1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.620 2.300 2.740 ;
        RECT  2.080 2.460 2.300 2.740 ;
        RECT  1.460 0.620 2.300 0.820 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.280 0.700 1.560 ;
        RECT  0.500 1.100 0.700 1.560 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.100 1.960 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.020 -0.280 2.300 0.420 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.330 -0.280 0.610 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.670 2.800 1.310 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.440 2.480 1.880 2.640 ;
        RECT  1.660 0.980 1.880 2.640 ;
        RECT  0.440 2.120 0.600 2.640 ;
        RECT  0.340 2.120 0.600 2.400 ;
        RECT  1.140 0.980 1.880 1.140 ;
        RECT  1.140 0.780 1.300 1.140 ;
        RECT  0.330 0.780 1.300 0.940 ;
    END
END AN2B1CHD

MACRO AN2B1EHD
    CLASS CORE ;
    FOREIGN AN2B1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.460 2.700 2.740 ;
        RECT  2.480 2.460 2.700 2.740 ;
        RECT  2.480 0.460 2.700 0.740 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.320 1.900 1.960 ;
        RECT  1.650 1.520 1.900 1.800 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.680 0.700 1.960 ;
        RECT  0.500 1.440 0.700 1.960 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.440 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.330 -0.280 0.610 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.890 2.800 1.530 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.380 2.120 2.280 2.280 ;
        RECT  2.120 0.700 2.280 2.280 ;
        RECT  2.080 1.400 2.300 1.680 ;
        RECT  0.930 0.700 2.280 0.860 ;
        RECT  0.300 2.240 1.080 2.400 ;
        RECT  0.920 1.020 1.080 2.400 ;
        RECT  0.300 2.180 0.580 2.400 ;
        RECT  0.450 1.020 1.080 1.180 ;
        RECT  0.450 0.780 0.610 1.180 ;
        RECT  0.330 0.780 0.610 0.940 ;
    END
END AN2B1EHD

MACRO AN2B1HHD
    CLASS CORE ;
    FOREIGN AN2B1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.460 2.700 2.740 ;
        RECT  2.500 2.460 2.760 2.740 ;
        RECT  2.440 0.460 2.700 0.740 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.320 1.900 1.960 ;
        RECT  1.650 1.520 1.900 1.800 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.680 0.700 1.960 ;
        RECT  0.500 1.440 0.700 1.960 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.810 -0.280 2.090 0.440 ;
        RECT  3.140 -0.280 3.420 0.780 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.330 -0.280 0.610 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.980 2.800 2.260 3.480 ;
        RECT  3.100 2.800 3.380 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.760 2.800 1.040 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.380 2.120 2.280 2.280 ;
        RECT  2.120 0.700 2.280 2.280 ;
        RECT  2.080 1.400 2.300 1.680 ;
        RECT  0.930 0.700 2.280 0.860 ;
        RECT  0.300 2.240 1.080 2.400 ;
        RECT  0.920 1.020 1.080 2.400 ;
        RECT  0.300 2.180 0.580 2.400 ;
        RECT  0.450 1.020 1.080 1.180 ;
        RECT  0.450 0.780 0.610 1.180 ;
        RECT  0.330 0.780 0.610 0.940 ;
    END
END AN2B1HHD

MACRO AN2B1KHD
    CLASS CORE ;
    FOREIGN AN2B1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.360 0.640 5.780 0.840 ;
        RECT  4.360 2.100 5.780 2.300 ;
        RECT  4.900 0.640 5.100 2.300 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.780 1.680 ;
        RECT  2.500 1.240 2.700 1.880 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.100 0.700 1.660 ;
        RECT  0.400 1.280 0.700 1.560 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.790 -0.280 3.070 0.420 ;
        RECT  3.840 -0.280 4.120 0.580 ;
        RECT  4.940 -0.280 5.220 0.420 ;
        RECT  6.020 -0.280 6.300 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.110 -0.280 0.390 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 2.800 1.320 3.480 ;
        RECT  2.280 2.560 2.560 3.480 ;
        RECT  3.740 2.100 3.900 3.480 ;
        RECT  4.940 2.560 5.220 3.480 ;
        RECT  6.020 2.560 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.660 2.120 3.480 2.280 ;
        RECT  3.320 0.920 3.480 2.280 ;
        RECT  3.320 1.460 4.500 1.620 ;
        RECT  1.660 0.920 3.480 1.080 ;
        RECT  1.240 0.600 1.400 0.920 ;
        RECT  1.240 0.600 3.640 0.760 ;
        RECT  0.880 0.520 1.080 2.280 ;
        RECT  0.740 1.840 1.080 2.120 ;
        RECT  0.740 0.640 1.080 0.920 ;
    END
END AN2B1KHD

MACRO AN2CHD
    CLASS CORE ;
    FOREIGN AN2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.720 1.900 2.440 ;
        RECT  1.680 2.160 1.900 2.440 ;
        RECT  1.680 0.720 1.900 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.680 1.100 1.960 ;
        RECT  0.900 1.320 1.100 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.280 0.700 1.560 ;
        RECT  0.500 1.100 0.700 1.560 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  1.050 -0.280 1.330 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.320 2.800 1.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.540 2.120 1.460 2.280 ;
        RECT  1.300 0.740 1.460 2.280 ;
        RECT  1.300 1.400 1.500 1.680 ;
        RECT  0.120 0.740 1.460 0.900 ;
    END
END AN2CHD

MACRO AN2EHD
    CLASS CORE ;
    FOREIGN AN2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.460 1.900 2.740 ;
        RECT  1.680 2.460 1.900 2.740 ;
        RECT  1.680 0.460 1.900 0.740 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.100 1.960 ;
        RECT  0.860 1.570 1.100 1.850 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.280 0.700 1.560 ;
        RECT  0.500 1.060 0.700 1.560 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  1.050 -0.280 1.330 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.320 2.800 0.600 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.540 2.120 1.460 2.280 ;
        RECT  1.300 0.700 1.460 2.280 ;
        RECT  1.300 1.400 1.500 1.680 ;
        RECT  0.120 0.700 1.460 0.860 ;
    END
END AN2EHD

MACRO AN2HHD
    CLASS CORE ;
    FOREIGN AN2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.460 0.440 2.300 0.640 ;
        RECT  2.100 0.440 2.300 2.300 ;
        RECT  1.760 2.100 2.300 2.300 ;
        RECT  1.760 2.100 1.920 2.380 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.320 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.480 -0.280 2.640 0.920 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.940 -0.280 1.220 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.620 1.460 3.480 ;
        RECT  2.260 2.800 2.540 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.160 2.300 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 2.240 1.520 2.400 ;
        RECT  1.360 0.800 1.520 2.400 ;
        RECT  1.360 1.400 1.600 1.680 ;
        RECT  0.520 0.800 1.520 0.960 ;
        RECT  0.520 0.480 0.680 0.960 ;
        RECT  0.100 0.480 0.680 0.640 ;
        RECT  0.100 0.440 0.380 0.640 ;
    END
END AN2HHD

MACRO AN2KHD
    CLASS CORE ;
    FOREIGN AN2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.440 3.100 2.380 ;
        RECT  2.900 1.300 3.900 1.500 ;
        RECT  3.700 0.440 3.900 2.400 ;
        RECT  3.700 2.200 4.160 2.400 ;
        RECT  3.960 2.200 4.160 2.760 ;
        RECT  3.700 0.440 4.180 0.640 ;
        RECT  2.620 0.440 3.100 0.640 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.320 2.300 1.960 ;
        RECT  2.020 1.400 2.300 1.680 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.080 1.360 1.500 1.560 ;
        RECT  1.300 0.920 1.500 1.560 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.300 -0.280 3.460 0.680 ;
        RECT  4.420 -0.280 4.700 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  2.100 -0.280 2.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 2.580 1.500 3.480 ;
        RECT  2.340 2.620 2.620 3.480 ;
        RECT  3.380 2.620 3.660 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 2.120 2.740 2.280 ;
        RECT  2.580 0.800 2.740 2.280 ;
        RECT  1.760 0.800 2.740 0.960 ;
        RECT  1.760 0.520 1.920 0.960 ;
        RECT  0.130 0.520 1.920 0.680 ;
    END
END AN2KHD

MACRO AN3B1CHD
    CLASS CORE ;
    FOREIGN AN3B1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.720 3.900 2.440 ;
        RECT  3.680 2.160 3.900 2.440 ;
        RECT  3.680 0.720 3.900 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.840 1.680 3.100 1.960 ;
        RECT  2.900 1.400 3.100 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.460 1.520 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.100 0.700 1.660 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.050 -0.280 3.330 0.440 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.250 -0.280 0.530 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.560 2.140 3.480 ;
        RECT  3.030 2.560 3.310 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.240 2.800 0.520 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.300 2.180 1.580 2.440 ;
        RECT  1.300 2.180 3.480 2.340 ;
        RECT  3.280 0.600 3.480 2.340 ;
        RECT  1.540 0.600 3.480 0.760 ;
        RECT  0.880 2.060 1.100 2.340 ;
        RECT  0.900 0.640 1.100 2.340 ;
        RECT  0.900 1.680 1.180 1.960 ;
        RECT  0.880 0.640 1.100 0.920 ;
    END
END AN3B1CHD

MACRO AN3B1EHD
    CLASS CORE ;
    FOREIGN AN3B1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.460 3.900 2.740 ;
        RECT  3.680 2.460 3.900 2.740 ;
        RECT  3.680 0.460 3.900 0.740 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.400 3.100 1.960 ;
        RECT  2.840 1.620 3.100 1.900 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.350 2.460 1.630 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.100 0.700 1.660 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.050 -0.280 3.330 0.440 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.250 -0.280 0.530 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.560 2.140 3.480 ;
        RECT  3.030 2.560 3.310 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.240 2.800 0.520 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.300 2.120 1.580 2.400 ;
        RECT  1.300 2.180 3.480 2.340 ;
        RECT  3.280 0.600 3.480 2.340 ;
        RECT  1.540 0.600 3.480 0.760 ;
        RECT  0.880 2.060 1.100 2.340 ;
        RECT  0.900 0.640 1.100 2.340 ;
        RECT  0.900 1.620 1.180 1.900 ;
        RECT  0.880 0.640 1.100 0.920 ;
    END
END AN3B1EHD

MACRO AN3B1HHD
    CLASS CORE ;
    FOREIGN AN3B1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.460 3.900 2.740 ;
        RECT  3.540 2.460 3.900 2.740 ;
        RECT  3.540 0.460 3.900 0.740 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.580 2.860 1.860 ;
        RECT  2.500 1.400 2.700 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.350 2.320 1.630 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.100 0.700 1.660 ;
        RECT  0.400 1.280 0.700 1.560 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.910 -0.280 3.190 0.440 ;
        RECT  4.240 -0.280 4.520 0.640 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.110 -0.280 0.390 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.720 2.800 2.000 3.480 ;
        RECT  2.890 2.800 3.170 3.480 ;
        RECT  4.240 2.580 4.520 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.220 2.480 1.480 2.760 ;
        RECT  1.220 2.480 3.340 2.640 ;
        RECT  3.180 0.600 3.340 2.640 ;
        RECT  3.180 1.400 3.360 1.680 ;
        RECT  1.400 0.600 3.340 0.760 ;
        RECT  0.740 2.060 1.100 2.340 ;
        RECT  0.900 0.640 1.100 2.340 ;
        RECT  0.740 0.640 1.100 0.920 ;
    END
END AN3B1HHD

MACRO AN3B2BHD
    CLASS CORE ;
    FOREIGN AN3B2BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.620 3.100 2.740 ;
        RECT  2.870 2.460 3.100 2.740 ;
        RECT  1.650 0.620 3.100 0.820 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.390 1.280 0.700 1.560 ;
        RECT  0.500 1.100 0.700 1.560 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.320 1.500 1.960 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.320 2.300 2.370 ;
        RECT  2.030 1.400 2.300 1.680 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.930 -0.280 1.210 0.420 ;
        RECT  2.250 -0.280 2.530 0.420 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.330 -0.280 0.610 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.670 2.800 0.950 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.110 2.600 2.690 2.760 ;
        RECT  2.530 0.980 2.690 2.760 ;
        RECT  0.420 2.480 1.270 2.640 ;
        RECT  0.420 2.120 0.580 2.640 ;
        RECT  0.360 2.120 0.580 2.400 ;
        RECT  1.330 0.980 2.690 1.140 ;
        RECT  1.330 0.780 1.490 1.140 ;
        RECT  0.330 0.780 1.490 0.940 ;
    END
END AN3B2BHD

MACRO AN3B2EHD
    CLASS CORE ;
    FOREIGN AN3B2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.460 4.300 2.740 ;
        RECT  4.080 2.460 4.300 2.740 ;
        RECT  4.080 0.460 4.300 0.740 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.320 3.500 1.960 ;
        RECT  3.240 1.620 3.500 1.900 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.320 0.700 1.960 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.350 1.160 1.630 ;
        RECT  0.900 0.920 1.100 1.630 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.450 -0.280 3.730 0.440 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.260 2.560 2.540 3.480 ;
        RECT  3.430 2.560 3.710 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.180 3.880 2.340 ;
        RECT  3.660 0.600 3.880 2.340 ;
        RECT  2.000 0.600 2.220 0.880 ;
        RECT  2.000 0.600 3.880 0.760 ;
        RECT  0.120 2.060 0.320 2.340 ;
        RECT  0.120 0.580 0.280 2.340 ;
        RECT  2.640 1.360 2.920 1.570 ;
        RECT  1.660 1.360 2.920 1.520 ;
        RECT  1.660 0.580 1.820 1.520 ;
        RECT  0.120 0.960 0.320 1.240 ;
        RECT  0.120 0.580 1.820 0.740 ;
        RECT  1.280 2.060 1.480 2.340 ;
        RECT  1.320 0.960 1.480 2.340 ;
        RECT  1.320 1.680 2.160 1.840 ;
        RECT  1.280 0.960 1.480 1.240 ;
    END
END AN3B2EHD

MACRO AN3B2HHD
    CLASS CORE ;
    FOREIGN AN3B2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.460 4.300 2.740 ;
        RECT  4.020 2.460 4.300 2.740 ;
        RECT  4.020 0.460 4.300 0.740 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.320 3.500 1.960 ;
        RECT  3.240 1.520 3.500 1.800 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.400 0.700 1.960 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.350 1.160 1.630 ;
        RECT  0.900 0.920 1.100 1.630 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.400 -0.280 3.680 0.420 ;
        RECT  4.740 -0.280 5.020 0.780 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.260 2.560 2.540 3.480 ;
        RECT  3.400 2.560 3.680 3.480 ;
        RECT  4.740 2.420 5.020 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.180 3.840 2.340 ;
        RECT  3.680 0.600 3.840 2.340 ;
        RECT  3.680 1.400 3.880 1.680 ;
        RECT  2.000 0.600 2.200 0.880 ;
        RECT  2.000 0.600 3.840 0.760 ;
        RECT  0.120 2.060 0.320 2.340 ;
        RECT  0.120 0.580 0.280 2.340 ;
        RECT  2.640 1.260 2.920 1.560 ;
        RECT  1.660 1.260 2.920 1.420 ;
        RECT  1.660 0.580 1.820 1.420 ;
        RECT  0.120 0.960 0.320 1.240 ;
        RECT  0.120 0.580 1.820 0.740 ;
        RECT  1.280 2.060 1.480 2.340 ;
        RECT  1.320 0.960 1.480 2.340 ;
        RECT  1.320 1.580 2.160 1.740 ;
        RECT  1.280 0.960 1.480 1.240 ;
    END
END AN3B2HHD

MACRO AN3CHD
    CLASS CORE ;
    FOREIGN AN3CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.720 2.700 2.440 ;
        RECT  2.480 2.160 2.700 2.440 ;
        RECT  2.480 0.720 2.700 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.260 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.640 0.740 2.020 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.680 1.900 1.960 ;
        RECT  1.700 1.320 1.900 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  1.850 -0.280 2.130 0.440 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.830 2.560 2.110 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.180 0.380 2.400 ;
        RECT  0.100 2.180 2.280 2.340 ;
        RECT  2.060 0.600 2.280 2.340 ;
        RECT  0.340 0.600 2.280 0.760 ;
    END
END AN3CHD

MACRO AN3EHD
    CLASS CORE ;
    FOREIGN AN3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.440 2.700 2.760 ;
        RECT  2.480 2.480 2.700 2.760 ;
        RECT  2.480 0.440 2.700 0.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.680 1.260 1.960 ;
        RECT  0.900 1.320 1.100 2.020 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.880 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.680 1.900 1.960 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  1.850 -0.280 2.130 0.440 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.830 2.560 2.110 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.180 0.380 2.400 ;
        RECT  0.100 2.180 2.280 2.340 ;
        RECT  2.120 0.600 2.280 2.340 ;
        RECT  2.100 1.400 2.300 1.680 ;
        RECT  0.340 0.600 2.280 0.760 ;
    END
END AN3EHD

MACRO AN3HHD
    CLASS CORE ;
    FOREIGN AN3HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.440 2.700 2.760 ;
        RECT  2.480 2.480 2.700 2.760 ;
        RECT  2.480 0.440 2.700 0.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.660 1.120 1.940 ;
        RECT  0.900 1.560 1.100 2.080 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.400 0.380 1.680 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.890 ;
        RECT  1.640 1.340 1.900 1.620 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.010 -0.280 3.290 0.660 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  1.640 -0.280 1.920 0.660 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.830 2.560 2.110 3.480 ;
        RECT  3.010 2.560 3.290 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.670 2.560 0.950 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.240 0.380 2.460 ;
        RECT  0.100 2.240 2.280 2.400 ;
        RECT  2.120 0.820 2.280 2.400 ;
        RECT  2.100 1.400 2.300 1.680 ;
        RECT  1.320 0.820 2.280 0.980 ;
        RECT  1.320 0.520 1.480 0.980 ;
        RECT  0.100 0.520 0.380 0.740 ;
        RECT  0.100 0.520 1.480 0.680 ;
    END
END AN3HHD

MACRO AN4B1BHD
    CLASS CORE ;
    FOREIGN AN4B1BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.790 3.500 2.640 ;
        RECT  3.280 2.360 3.500 2.640 ;
        RECT  2.660 0.790 3.500 0.990 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.260 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.640 0.740 2.020 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.880 ;
        RECT  2.380 1.240 2.700 1.520 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.680 1.900 1.960 ;
        RECT  1.700 1.320 1.900 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.220 -0.280 3.500 0.420 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  1.850 -0.280 2.130 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.830 2.560 2.110 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.180 0.380 2.400 ;
        RECT  0.100 2.180 3.060 2.340 ;
        RECT  2.900 1.240 3.060 2.340 ;
        RECT  2.060 0.600 2.220 2.340 ;
        RECT  0.340 0.600 2.220 0.760 ;
    END
END AN4B1BHD

MACRO AN4B1EHD
    CLASS CORE ;
    FOREIGN AN4B1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.000 0.440 3.200 0.990 ;
        RECT  3.300 0.790 3.500 2.360 ;
        RECT  3.000 0.790 4.140 0.990 ;
        RECT  2.590 0.440 3.200 0.640 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.260 1.620 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.640 0.740 2.020 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 1.240 2.700 1.880 ;
        RECT  4.120 1.240 4.280 2.680 ;
        RECT  2.380 2.520 4.280 2.680 ;
        RECT  2.380 1.240 2.540 2.680 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.640 1.680 1.900 1.960 ;
        RECT  1.700 1.320 1.900 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.360 -0.280 3.520 0.480 ;
        RECT  4.420 -0.280 4.700 0.420 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  1.850 -0.280 2.130 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.830 2.560 2.110 3.480 ;
        RECT  4.420 2.780 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.180 0.380 2.400 ;
        RECT  0.100 2.180 2.220 2.340 ;
        RECT  2.060 0.600 2.220 2.340 ;
        RECT  2.060 0.920 2.840 1.080 ;
        RECT  0.340 0.600 2.220 0.760 ;
    END
END AN4B1EHD

MACRO AN4B1HHD
    CLASS CORE ;
    FOREIGN AN4B1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.460 0.600 4.890 0.800 ;
        RECT  4.690 0.440 5.540 0.640 ;
        RECT  5.340 0.440 5.540 0.990 ;
        RECT  5.700 0.790 5.900 2.360 ;
        RECT  5.340 0.790 6.540 0.990 ;
        RECT  3.020 0.600 3.220 2.360 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.260 1.620 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.620 0.740 2.020 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.380 1.520 3.540 2.680 ;
        RECT  2.380 2.520 3.540 2.680 ;
        RECT  4.500 1.520 4.700 2.280 ;
        RECT  3.380 1.520 5.480 1.680 ;
        RECT  5.320 1.520 5.480 2.680 ;
        RECT  6.520 1.240 6.680 2.680 ;
        RECT  5.320 2.520 6.680 2.680 ;
        RECT  2.380 1.460 2.540 2.680 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.320 1.900 1.960 ;
        RECT  1.640 1.540 1.900 1.820 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.020 -0.280 3.300 0.420 ;
        RECT  4.140 -0.280 4.420 0.420 ;
        RECT  5.700 -0.280 5.980 0.420 ;
        RECT  6.820 -0.280 7.100 0.420 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  1.850 -0.280 2.130 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.830 2.560 2.110 3.480 ;
        RECT  3.940 2.580 4.970 3.480 ;
        RECT  6.820 2.780 7.100 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.660 2.560 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.020 0.980 5.180 1.260 ;
        RECT  3.400 1.040 5.180 1.200 ;
        RECT  0.100 2.180 0.380 2.400 ;
        RECT  0.100 2.180 2.220 2.340 ;
        RECT  2.060 0.600 2.220 2.340 ;
        RECT  2.560 1.040 2.840 1.260 ;
        RECT  2.060 1.040 2.840 1.200 ;
        RECT  0.340 0.600 2.220 0.760 ;
    END
END AN4B1HHD

MACRO AN4CHD
    CLASS CORE ;
    FOREIGN AN4CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.720 2.300 2.760 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.680 1.100 1.960 ;
        RECT  0.900 1.320 1.100 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.360 1.280 0.700 1.560 ;
        RECT  0.500 1.100 0.700 1.560 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.680 3.160 1.960 ;
        RECT  2.900 1.400 3.100 1.960 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.280 3.640 1.560 ;
        RECT  3.300 1.100 3.500 1.560 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.670 -0.280 2.950 0.460 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  1.050 -0.280 1.330 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.040 2.800 3.680 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.320 2.800 1.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.520 2.120 3.460 2.280 ;
        RECT  2.520 0.740 2.680 2.280 ;
        RECT  2.520 0.740 3.880 0.900 ;
        RECT  0.540 2.120 1.480 2.280 ;
        RECT  1.320 0.740 1.480 2.280 ;
        RECT  1.300 1.400 1.500 1.680 ;
        RECT  0.120 0.740 1.480 0.900 ;
    END
END AN4CHD

MACRO AN4EHD
    CLASS CORE ;
    FOREIGN AN4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 2.100 2.220 2.300 ;
        RECT  1.700 0.440 1.900 2.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.680 1.100 1.960 ;
        RECT  0.900 1.320 1.100 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.120 1.360 0.700 1.560 ;
        RECT  0.500 1.100 0.700 1.560 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.840 3.500 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.400 4.040 1.680 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 -0.280 2.620 0.440 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  1.050 -0.280 1.330 0.440 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.440 2.800 4.080 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.320 2.800 1.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.980 2.020 3.860 2.180 ;
        RECT  2.980 0.440 3.140 2.180 ;
        RECT  2.120 0.920 2.280 1.660 ;
        RECT  2.120 0.920 3.140 1.080 ;
        RECT  4.000 0.440 4.280 0.660 ;
        RECT  2.980 0.440 4.280 0.600 ;
        RECT  1.320 2.520 2.680 2.680 ;
        RECT  2.520 1.460 2.680 2.680 ;
        RECT  1.320 0.740 1.480 2.680 ;
        RECT  0.540 2.120 1.480 2.280 ;
        RECT  2.520 1.460 2.820 1.740 ;
        RECT  0.120 0.740 1.480 0.900 ;
    END
END AN4EHD

MACRO AN4HHD
    CLASS CORE ;
    FOREIGN AN4HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.960 3.100 2.300 ;
        RECT  1.940 2.100 3.100 2.300 ;
        RECT  2.900 0.960 3.900 1.160 ;
        RECT  3.700 0.960 3.900 2.300 ;
        RECT  3.700 2.100 4.220 2.300 ;
        RECT  1.940 0.440 2.140 2.300 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.120 1.380 0.700 1.580 ;
        RECT  0.500 1.100 0.700 1.580 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.840 5.500 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.400 6.040 1.680 ;
        RECT  5.700 1.240 5.900 1.760 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.500 -0.280 2.780 0.440 ;
        RECT  4.340 -0.280 4.620 0.440 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  1.160 -0.280 1.440 0.440 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.200 2.800 1.380 3.480 ;
        RECT  3.060 2.800 3.340 3.480 ;
        RECT  5.080 2.360 5.240 3.480 ;
        RECT  5.080 2.800 6.200 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  1.100 2.420 1.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.980 2.020 5.860 2.180 ;
        RECT  4.980 0.440 5.140 2.180 ;
        RECT  4.120 0.600 4.280 1.660 ;
        RECT  2.360 0.600 2.520 1.660 ;
        RECT  2.360 0.600 5.140 0.760 ;
        RECT  6.000 0.440 6.280 0.660 ;
        RECT  4.980 0.440 6.280 0.600 ;
        RECT  1.560 2.480 4.790 2.640 ;
        RECT  4.630 1.360 4.790 2.640 ;
        RECT  3.320 1.420 3.480 2.640 ;
        RECT  1.560 0.600 1.720 2.640 ;
        RECT  0.500 2.100 1.720 2.260 ;
        RECT  4.630 1.460 4.820 1.740 ;
        RECT  0.120 0.600 1.720 0.760 ;
    END
END AN4HHD

MACRO ANTHD
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 0.540 0.580 1.160 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 0.800 3.480 ;
        END
    END VCC
END ANTHD

MACRO AO112CHD
    CLASS CORE ;
    FOREIGN AO112CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.720 3.500 2.440 ;
        RECT  3.280 2.160 3.500 2.440 ;
        RECT  3.280 0.720 3.500 1.000 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.320 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.630 -0.280 2.930 0.460 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.140 2.460 0.420 2.680 ;
        RECT  0.140 2.460 0.880 2.620 ;
        RECT  0.720 2.160 0.880 2.620 ;
        RECT  0.860 0.740 1.020 2.320 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AO112CHD

MACRO AO112EHD
    CLASS CORE ;
    FOREIGN AO112EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  3.280 0.460 3.500 0.740 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.320 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.650 -0.280 2.930 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.880 2.540 ;
        RECT  0.720 2.060 0.880 2.540 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AO112EHD

MACRO AO112HHD
    CLASS CORE ;
    FOREIGN AO112HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  3.280 0.460 3.500 0.740 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.320 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.790 -0.280 4.070 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.780 2.800 4.060 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.680 2.540 ;
        RECT  0.520 1.980 0.680 2.540 ;
        RECT  0.520 1.980 1.020 2.140 ;
        RECT  0.860 0.740 1.020 2.140 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.020 2.480 2.420 2.640 ;
    END
END AO112HHD

MACRO AO112KHD
    CLASS CORE ;
    FOREIGN AO112KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  4.400 0.460 4.700 0.740 ;
        RECT  3.300 1.300 4.700 1.500 ;
        RECT  4.500 0.460 4.700 2.740 ;
        RECT  4.400 2.460 4.700 2.740 ;
        RECT  3.280 0.460 3.500 0.740 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.320 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.780 -0.280 4.060 0.400 ;
        RECT  5.100 -0.280 5.380 0.780 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.780 2.800 4.060 3.480 ;
        RECT  5.100 2.420 5.380 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.880 2.540 ;
        RECT  0.720 2.060 0.880 2.540 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AO112KHD

MACRO AO12CHD
    CLASS CORE ;
    FOREIGN AO12CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.460 2.700 2.340 ;
        RECT  2.480 2.060 2.700 2.340 ;
        RECT  2.480 0.460 2.700 0.740 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.320 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.880 ;
        RECT  1.640 1.400 1.900 1.680 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.980 -0.280 1.260 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.820 2.800 2.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.580 2.280 2.280 2.440 ;
        RECT  2.120 0.780 2.280 2.440 ;
        RECT  1.520 0.780 1.800 1.020 ;
        RECT  0.100 0.780 2.280 0.940 ;
        RECT  0.100 0.720 0.380 0.940 ;
        RECT  0.100 2.600 1.500 2.760 ;
        RECT  0.100 2.540 0.380 2.760 ;
    END
END AO12CHD

MACRO AO12EHD
    CLASS CORE ;
    FOREIGN AO12EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.460 2.700 2.740 ;
        RECT  2.480 2.460 2.700 2.740 ;
        RECT  2.480 0.460 2.700 0.740 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.320 1.100 1.960 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.040 0.700 1.560 ;
        RECT  0.340 1.260 0.700 1.540 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.880 ;
        RECT  1.640 1.340 1.900 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  1.140 -0.280 1.420 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.860 2.800 2.140 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.740 2.280 2.280 2.440 ;
        RECT  2.120 0.780 2.280 2.440 ;
        RECT  1.520 0.780 1.800 0.960 ;
        RECT  1.520 0.780 2.280 0.940 ;
        RECT  1.520 0.560 1.680 0.960 ;
        RECT  0.100 0.560 1.680 0.720 ;
        RECT  0.100 0.500 0.380 0.720 ;
        RECT  0.220 2.600 1.580 2.760 ;
        RECT  0.100 2.380 0.380 2.700 ;
    END
END AO12EHD

MACRO AO12HHD
    CLASS CORE ;
    FOREIGN AO12HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.440 2.450 2.700 2.730 ;
        RECT  2.500 0.460 2.740 0.740 ;
        RECT  2.500 0.460 2.700 2.730 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.320 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.880 ;
        RECT  1.640 1.400 1.900 1.680 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.960 -0.280 2.240 0.400 ;
        RECT  3.140 -0.280 3.420 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.980 -0.280 1.260 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.140 2.420 3.420 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.740 2.800 2.020 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.580 2.480 2.280 2.640 ;
        RECT  2.120 0.780 2.280 2.640 ;
        RECT  2.100 1.400 2.300 1.680 ;
        RECT  1.520 0.780 1.800 1.020 ;
        RECT  0.100 0.780 2.280 0.940 ;
        RECT  0.100 0.720 0.380 0.940 ;
        RECT  0.100 2.140 0.380 2.360 ;
        RECT  0.100 2.140 1.460 2.300 ;
    END
END AO12HHD

MACRO AO12KHD
    CLASS CORE ;
    FOREIGN AO12KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.440 2.450 2.700 2.730 ;
        RECT  2.500 0.460 2.800 0.740 ;
        RECT  2.500 1.700 3.900 1.900 ;
        RECT  3.700 0.460 3.900 2.670 ;
        RECT  3.700 0.460 3.920 0.740 ;
        RECT  3.700 2.510 4.180 2.670 ;
        RECT  2.500 0.460 2.700 2.730 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.780 ;
        RECT  1.640 1.400 1.900 1.680 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.020 -0.280 2.300 0.400 ;
        RECT  3.140 -0.280 3.420 0.400 ;
        RECT  4.260 -0.280 4.540 0.400 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.980 -0.280 1.260 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.140 2.420 3.420 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  1.740 2.800 2.020 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 2.480 2.280 2.640 ;
        RECT  2.120 0.780 2.280 2.640 ;
        RECT  0.100 0.780 2.280 0.940 ;
        RECT  0.100 0.720 0.380 0.940 ;
        RECT  0.100 2.080 0.380 2.360 ;
        RECT  0.100 2.140 1.460 2.300 ;
    END
END AO12KHD

MACRO AO13CHD
    CLASS CORE ;
    FOREIGN AO13CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.720 3.500 2.440 ;
        RECT  3.280 2.160 3.500 2.440 ;
        RECT  3.280 0.720 3.500 1.000 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.380 2.580 ;
        RECT  0.100 2.380 0.800 2.540 ;
        RECT  0.640 2.000 0.800 2.540 ;
        RECT  0.640 2.000 1.020 2.160 ;
        RECT  0.860 0.740 1.020 2.160 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.420 2.380 2.580 ;
    END
END AO13CHD

MACRO AO13EHD
    CLASS CORE ;
    FOREIGN AO13EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  3.280 0.460 3.500 0.740 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.800 2.540 ;
        RECT  0.640 2.060 0.800 2.540 ;
        RECT  0.640 2.060 1.020 2.220 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AO13EHD

MACRO AO13HHD
    CLASS CORE ;
    FOREIGN AO13HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  3.280 0.460 3.500 0.740 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.780 -0.280 4.060 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.780 2.800 4.060 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.800 2.540 ;
        RECT  0.640 2.060 0.800 2.540 ;
        RECT  0.640 2.060 1.020 2.220 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AO13HHD

MACRO AO13KHD
    CLASS CORE ;
    FOREIGN AO13KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  4.400 0.460 4.700 0.740 ;
        RECT  3.300 1.300 4.700 1.500 ;
        RECT  4.500 0.460 4.700 2.740 ;
        RECT  4.400 2.460 4.700 2.740 ;
        RECT  3.280 0.460 3.500 0.740 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.780 -0.280 4.060 0.400 ;
        RECT  5.100 -0.280 5.380 0.780 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.780 2.800 4.060 3.480 ;
        RECT  5.100 2.420 5.380 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.480 0.800 2.640 ;
        RECT  0.640 2.060 0.800 2.640 ;
        RECT  0.640 2.060 1.020 2.220 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AO13KHD

MACRO AO2222BHD
    CLASS CORE ;
    FOREIGN AO2222BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.560 6.300 2.280 ;
        RECT  5.510 2.080 6.300 2.280 ;
        RECT  5.020 0.560 6.300 0.760 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.900 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.900 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.900 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        RECT  3.260 1.340 3.500 1.620 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  6.020 -0.280 6.300 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.910 2.800 5.190 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.720 2.600 4.740 2.760 ;
        RECT  4.580 2.300 4.740 2.760 ;
        RECT  2.720 2.120 2.880 2.760 ;
        RECT  4.580 2.300 5.350 2.460 ;
        RECT  5.190 1.740 5.350 2.460 ;
        RECT  1.100 2.120 2.880 2.280 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.190 1.740 5.900 1.900 ;
        RECT  5.740 1.460 5.900 1.900 ;
        RECT  0.620 0.920 1.880 1.080 ;
        RECT  3.540 1.960 5.020 2.120 ;
        RECT  4.860 0.920 5.020 2.120 ;
        RECT  4.860 1.400 5.480 1.560 ;
        RECT  3.060 0.920 5.020 1.080 ;
        RECT  2.600 0.600 2.760 1.020 ;
        RECT  2.600 0.600 4.820 0.760 ;
        RECT  3.060 2.280 4.420 2.440 ;
        RECT  3.060 2.220 3.340 2.440 ;
        RECT  2.120 0.600 2.280 1.020 ;
        RECT  0.160 0.600 0.320 1.020 ;
        RECT  0.160 0.600 2.280 0.760 ;
        RECT  0.580 2.440 1.980 2.600 ;
    END
END AO2222BHD

MACRO AO2222CHD
    CLASS CORE ;
    FOREIGN AO2222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.560 6.300 2.300 ;
        RECT  5.510 2.100 6.300 2.300 ;
        RECT  5.020 0.560 6.300 0.760 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.900 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.900 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        RECT  3.260 1.340 3.500 1.620 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  6.020 -0.280 6.300 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.900 2.800 5.180 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.680 2.600 4.740 2.760 ;
        RECT  4.580 2.300 4.740 2.760 ;
        RECT  2.680 2.120 2.840 2.760 ;
        RECT  4.580 2.300 5.350 2.460 ;
        RECT  5.190 1.740 5.350 2.460 ;
        RECT  1.100 2.120 2.840 2.280 ;
        RECT  1.720 0.880 1.880 2.280 ;
        RECT  5.190 1.740 5.900 1.900 ;
        RECT  5.740 1.460 5.900 1.900 ;
        RECT  0.620 0.880 1.880 1.040 ;
        RECT  3.540 1.960 5.020 2.120 ;
        RECT  4.860 0.920 5.020 2.120 ;
        RECT  4.860 1.400 5.480 1.560 ;
        RECT  3.020 0.920 5.020 1.080 ;
        RECT  2.600 0.600 2.760 0.920 ;
        RECT  2.600 0.600 4.820 0.760 ;
        RECT  3.020 2.280 4.420 2.440 ;
        RECT  2.120 0.560 2.280 0.920 ;
        RECT  0.160 0.560 0.320 0.920 ;
        RECT  0.160 0.560 2.280 0.720 ;
        RECT  0.620 2.440 1.940 2.600 ;
    END
END AO2222CHD

MACRO AO2222EHD
    CLASS CORE ;
    FOREIGN AO2222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 0.600 7.900 2.280 ;
        RECT  5.360 2.120 7.900 2.280 ;
        RECT  5.900 0.600 7.900 0.760 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.900 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.900 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.370 4.740 1.650 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  5.020 -0.280 5.300 0.760 ;
        RECT  7.500 -0.280 7.780 0.400 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.720 2.740 4.880 3.480 ;
        RECT  5.960 2.800 6.240 3.480 ;
        RECT  7.500 2.800 7.780 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.100 2.120 2.780 2.280 ;
        RECT  5.040 1.460 5.200 2.120 ;
        RECT  2.620 1.960 5.200 2.120 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.040 1.780 6.880 1.940 ;
        RECT  6.720 1.340 6.880 1.940 ;
        RECT  5.080 1.340 5.240 1.620 ;
        RECT  0.580 0.920 1.880 1.080 ;
        RECT  6.400 2.480 6.680 2.760 ;
        RECT  5.040 2.480 6.680 2.640 ;
        RECT  5.040 2.280 5.200 2.640 ;
        RECT  3.440 2.280 5.200 2.440 ;
        RECT  6.220 0.920 6.380 1.620 ;
        RECT  3.020 0.920 6.380 1.080 ;
        RECT  2.540 0.600 4.820 0.760 ;
        RECT  2.960 2.600 4.320 2.760 ;
        RECT  0.100 0.600 2.340 0.760 ;
        RECT  0.620 2.440 1.980 2.600 ;
    END
END AO2222EHD

MACRO AO2222HHD
    CLASS CORE ;
    FOREIGN AO2222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.600 9.500 2.280 ;
        RECT  5.320 2.120 9.500 2.280 ;
        RECT  5.860 0.600 9.500 0.760 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.900 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.900 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  5.020 -0.280 5.300 0.760 ;
        RECT  6.740 -0.280 7.020 0.400 ;
        RECT  9.220 -0.280 9.500 0.400 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.290 2.440 2.570 3.480 ;
        RECT  4.580 2.800 4.860 3.480 ;
        RECT  5.920 2.800 6.200 3.480 ;
        RECT  7.060 2.800 7.340 3.480 ;
        RECT  7.980 2.800 8.260 3.480 ;
        RECT  9.220 2.800 9.500 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.100 2.120 2.780 2.280 ;
        RECT  5.000 1.340 5.160 2.120 ;
        RECT  2.620 1.960 5.160 2.120 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.000 1.780 9.060 1.940 ;
        RECT  8.900 1.340 9.060 1.940 ;
        RECT  7.520 1.340 7.680 1.940 ;
        RECT  6.580 1.340 6.740 1.940 ;
        RECT  5.000 1.340 5.200 1.620 ;
        RECT  0.580 0.920 1.880 1.080 ;
        RECT  8.420 2.480 8.700 2.760 ;
        RECT  6.360 2.480 6.640 2.760 ;
        RECT  4.500 2.480 8.700 2.640 ;
        RECT  4.500 2.280 4.660 2.640 ;
        RECT  3.440 2.280 4.660 2.440 ;
        RECT  8.300 0.920 8.460 1.620 ;
        RECT  6.100 0.920 6.260 1.620 ;
        RECT  3.020 0.920 8.460 1.080 ;
        RECT  2.540 0.600 4.820 0.760 ;
        RECT  2.920 2.600 4.320 2.760 ;
        RECT  0.100 0.600 2.340 0.760 ;
        RECT  0.620 2.440 1.980 2.600 ;
    END
END AO2222HHD

MACRO AO222CHD
    CLASS CORE ;
    FOREIGN AO222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 0.920 4.700 2.280 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.250 1.100 1.880 ;
        RECT  0.860 1.370 1.100 1.650 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.340 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.580 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.540 1.650 ;
        RECT  1.300 1.250 1.500 1.880 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.250 2.300 1.770 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.280 3.990 0.400 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  1.020 -0.280 1.300 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.840 2.600 4.120 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  2.660 2.600 2.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.660 1.960 4.300 2.120 ;
        RECT  4.140 0.780 4.300 2.120 ;
        RECT  1.660 1.900 1.940 2.120 ;
        RECT  0.100 0.780 4.300 0.940 ;
        RECT  0.580 2.280 3.500 2.440 ;
        RECT  0.100 2.600 2.500 2.760 ;
        RECT  0.100 2.540 0.380 2.760 ;
    END
END AO222CHD

MACRO AO222EHD
    CLASS CORE ;
    FOREIGN AO222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 0.520 4.700 2.680 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.250 1.100 1.880 ;
        RECT  0.860 1.370 1.100 1.650 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.340 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.240 3.900 1.760 ;
        RECT  3.660 1.340 3.900 1.620 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.540 1.650 ;
        RECT  1.300 1.250 1.500 1.880 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.250 2.300 1.770 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.280 3.990 0.400 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  1.020 -0.280 1.300 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.860 2.620 4.140 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  2.780 2.620 3.060 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.660 1.840 1.880 2.120 ;
        RECT  1.720 0.700 1.880 2.120 ;
        RECT  4.140 0.700 4.300 1.660 ;
        RECT  0.100 0.700 4.300 0.860 ;
        RECT  0.580 2.280 2.200 2.440 ;
        RECT  2.040 2.060 2.200 2.440 ;
        RECT  2.040 2.060 3.620 2.220 ;
        RECT  0.100 2.600 2.600 2.760 ;
        RECT  2.360 2.380 2.600 2.760 ;
        RECT  0.100 2.540 0.380 2.760 ;
    END
END AO222EHD

MACRO AO222HHD
    CLASS CORE ;
    FOREIGN AO222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.300 0.900 5.100 1.100 ;
        RECT  4.900 0.900 5.100 2.300 ;
        RECT  4.310 2.100 5.100 2.300 ;
        RECT  4.300 2.100 5.100 2.260 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.760 ;
        RECT  1.540 1.370 1.900 1.650 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.620 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.860 1.370 1.100 1.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.360 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.690 -0.280 3.970 0.400 ;
        RECT  4.820 -0.280 5.100 0.600 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  1.260 -0.280 1.540 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 2.620 4.060 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  2.740 2.620 3.020 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.520 2.120 0.900 2.280 ;
        RECT  0.520 0.600 0.680 2.280 ;
        RECT  3.980 0.600 4.140 1.630 ;
        RECT  0.100 0.600 4.140 0.760 ;
        RECT  1.620 2.120 3.600 2.280 ;
        RECT  0.100 2.440 2.460 2.600 ;
    END
END AO222HHD

MACRO AO222KHD
    CLASS CORE ;
    FOREIGN AO222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.300 0.900 6.300 1.100 ;
        RECT  6.100 0.900 6.300 2.300 ;
        RECT  4.310 2.100 6.300 2.300 ;
        RECT  4.300 2.100 6.300 2.260 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.250 1.900 1.770 ;
        RECT  1.540 1.370 1.900 1.650 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.250 2.300 1.770 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.620 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.250 1.100 1.770 ;
        RECT  0.860 1.370 1.100 1.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.360 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.690 -0.280 3.970 0.400 ;
        RECT  4.820 -0.280 5.100 0.600 ;
        RECT  5.860 -0.280 6.140 0.600 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  1.260 -0.280 1.540 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 2.620 4.060 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  5.860 2.620 6.140 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  2.740 2.620 3.020 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.520 2.120 0.900 2.280 ;
        RECT  0.520 0.600 0.680 2.280 ;
        RECT  3.980 0.600 4.140 1.630 ;
        RECT  0.100 0.600 4.140 0.760 ;
        RECT  1.620 2.120 3.600 2.280 ;
        RECT  0.100 2.440 2.460 2.600 ;
    END
END AO222KHD

MACRO AO22CHD
    CLASS CORE ;
    FOREIGN AO22CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 0.920 3.500 2.280 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.140 1.620 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.760 ;
        RECT  2.480 1.390 2.700 1.670 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 1.940 1.620 ;
        RECT  1.700 1.240 1.900 1.760 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.640 -0.280 2.920 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 2.330 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.620 2.800 1.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 2.010 3.120 2.170 ;
        RECT  2.960 1.370 3.120 2.170 ;
        RECT  1.320 0.880 1.480 2.170 ;
        RECT  0.100 2.330 2.460 2.490 ;
    END
END AO22CHD

MACRO AO22EHD
    CLASS CORE ;
    FOREIGN AO22EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.680 0.520 3.900 2.680 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.140 1.620 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.880 1.390 3.100 1.670 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.340 2.340 1.620 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.040 -0.280 3.320 0.400 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  1.140 -0.280 1.420 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.480 3.380 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  2.020 2.800 2.300 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 2.160 3.520 2.320 ;
        RECT  3.360 0.560 3.520 2.320 ;
        RECT  0.560 0.920 0.720 2.320 ;
        RECT  0.100 0.920 0.720 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  2.060 0.560 3.520 0.720 ;
        RECT  0.100 2.480 2.860 2.640 ;
    END
END AO22EHD

MACRO AO22HHD
    CLASS CORE ;
    FOREIGN AO22HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.500 2.100 4.300 2.300 ;
        RECT  3.500 0.900 4.300 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.140 1.620 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.390 2.820 1.670 ;
        RECT  2.500 1.240 2.700 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 -0.280 3.200 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  1.260 -0.280 1.540 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  1.900 2.580 2.180 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 1.940 3.340 2.100 ;
        RECT  3.180 0.560 3.340 2.100 ;
        RECT  0.560 0.920 0.720 2.100 ;
        RECT  0.100 0.920 0.720 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.940 0.560 3.340 0.720 ;
        RECT  0.100 2.260 2.780 2.420 ;
    END
END AO22HHD

MACRO AO22KHD
    CLASS CORE ;
    FOREIGN AO22KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.900 5.500 2.300 ;
        RECT  3.500 2.100 5.500 2.300 ;
        RECT  3.500 0.900 5.500 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.140 1.620 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.390 2.820 1.670 ;
        RECT  2.500 1.240 2.700 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 -0.280 3.200 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  5.060 -0.280 5.340 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  1.260 -0.280 1.540 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  5.060 2.620 5.340 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  1.900 2.580 2.180 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 1.940 0.940 2.100 ;
        RECT  0.560 0.780 0.720 2.100 ;
        RECT  3.180 0.560 3.340 1.650 ;
        RECT  0.100 0.780 1.880 0.940 ;
        RECT  1.720 0.560 1.880 0.940 ;
        RECT  1.720 0.560 3.340 0.720 ;
        RECT  0.100 2.600 1.080 2.760 ;
        RECT  0.920 2.260 1.080 2.760 ;
        RECT  0.100 2.540 0.380 2.760 ;
        RECT  0.920 2.260 2.780 2.420 ;
    END
END AO22KHD

MACRO AOI112BHD
    CLASS CORE ;
    FOREIGN AOI112BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 2.380 0.880 2.540 ;
        RECT  0.860 0.700 1.020 2.220 ;
        RECT  0.100 0.700 3.100 0.900 ;
        RECT  2.900 0.700 3.100 2.600 ;
        RECT  0.720 2.060 0.880 2.540 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.650 -0.280 2.930 0.400 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AOI112BHD

MACRO AOI112EHD
    CLASS CORE ;
    FOREIGN AOI112EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.460 4.700 2.740 ;
        RECT  4.480 2.460 4.700 2.740 ;
        RECT  4.480 0.460 4.700 0.740 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.860 -0.280 4.140 0.400 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.860 2.800 4.140 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 1.840 3.500 2.120 ;
        RECT  3.300 0.960 3.500 2.120 ;
        RECT  3.300 1.400 4.300 1.680 ;
        RECT  3.280 0.960 3.500 1.240 ;
        RECT  0.100 2.380 0.880 2.540 ;
        RECT  0.720 2.060 0.880 2.540 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AOI112EHD

MACRO AOI112HHD
    CLASS CORE ;
    FOREIGN AOI112HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.460 4.700 2.740 ;
        RECT  4.340 2.460 4.700 2.740 ;
        RECT  4.340 0.460 4.700 0.740 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.700 -0.280 3.980 0.400 ;
        RECT  5.060 -0.280 5.340 0.780 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.700 2.800 3.980 3.480 ;
        RECT  5.060 2.420 5.340 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 1.840 3.500 2.120 ;
        RECT  3.300 0.960 3.500 2.120 ;
        RECT  3.300 1.400 4.140 1.680 ;
        RECT  3.280 0.960 3.500 1.240 ;
        RECT  0.100 2.380 0.880 2.540 ;
        RECT  0.720 2.060 0.880 2.540 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AOI112HHD

MACRO AOI112KHD
    CLASS CORE ;
    FOREIGN AOI112KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.460 4.700 2.740 ;
        RECT  4.340 2.460 4.700 2.740 ;
        RECT  4.500 1.400 5.900 1.680 ;
        RECT  5.700 0.460 5.900 2.740 ;
        RECT  5.700 0.460 6.060 0.740 ;
        RECT  5.700 2.460 6.060 2.740 ;
        RECT  4.340 0.460 4.700 0.740 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.280 1.500 1.560 ;
        RECT  1.300 1.060 1.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.280 2.020 1.560 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.700 -0.280 3.980 0.400 ;
        RECT  5.060 -0.280 5.340 0.780 ;
        RECT  6.420 -0.280 6.700 0.400 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.700 2.800 3.980 3.480 ;
        RECT  5.060 2.420 5.340 3.480 ;
        RECT  6.420 2.800 6.700 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 1.840 3.500 2.120 ;
        RECT  3.300 0.960 3.500 2.120 ;
        RECT  3.300 1.400 4.140 1.680 ;
        RECT  3.280 0.960 3.500 1.240 ;
        RECT  0.100 2.380 0.880 2.540 ;
        RECT  0.720 2.060 0.880 2.540 ;
        RECT  0.860 0.740 1.020 2.220 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  1.060 2.480 2.380 2.640 ;
    END
END AOI112KHD

MACRO AOI12CHD
    CLASS CORE ;
    FOREIGN AOI12CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.140 0.500 2.700 0.700 ;
        RECT  2.500 0.500 2.700 2.280 ;
        RECT  0.100 2.120 2.700 2.280 ;
        RECT  0.100 0.620 1.340 0.820 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.640 1.560 ;
        RECT  1.300 1.040 1.500 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.400 2.300 1.960 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.280 0.700 1.560 ;
        RECT  0.500 1.040 0.700 1.560 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 2.800 2.600 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.200 2.800 1.480 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.720 2.480 2.040 2.640 ;
    END
END AOI12CHD

MACRO AOI12EHD
    CLASS CORE ;
    FOREIGN AOI12EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.560 3.780 0.720 ;
        RECT  3.300 2.480 3.780 2.640 ;
        RECT  3.300 0.560 3.500 2.640 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.780 ;
        RECT  1.640 1.400 1.900 1.680 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  2.900 -0.280 3.180 0.400 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.980 -0.280 1.260 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.900 2.800 3.180 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  1.820 2.800 2.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.480 0.480 2.640 2.600 ;
        RECT  2.480 1.400 3.100 1.680 ;
        RECT  0.580 2.280 2.280 2.440 ;
        RECT  2.120 0.720 2.280 2.440 ;
        RECT  1.520 0.720 1.800 1.020 ;
        RECT  0.100 0.720 2.280 0.880 ;
        RECT  0.100 0.660 0.380 0.880 ;
        RECT  0.100 2.600 1.500 2.760 ;
        RECT  0.100 2.540 0.380 2.760 ;
    END
END AOI12EHD

MACRO AOI12HHD
    CLASS CORE ;
    FOREIGN AOI12HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.520 3.900 2.680 ;
        RECT  3.440 2.400 3.900 2.680 ;
        RECT  3.440 0.520 3.900 0.800 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.780 ;
        RECT  1.640 1.400 1.900 1.680 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.280 2.120 0.400 ;
        RECT  2.880 -0.280 3.160 0.400 ;
        RECT  4.200 -0.280 4.480 0.800 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.980 -0.280 1.260 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.880 2.800 3.160 3.480 ;
        RECT  4.200 2.420 4.480 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  1.740 2.800 2.020 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.440 0.960 2.640 2.120 ;
        RECT  2.440 1.400 2.760 1.680 ;
        RECT  0.620 2.480 2.280 2.640 ;
        RECT  2.120 0.780 2.280 2.640 ;
        RECT  1.460 0.780 1.740 1.020 ;
        RECT  0.100 0.780 2.280 0.940 ;
        RECT  0.100 0.720 0.380 0.940 ;
        RECT  0.100 2.080 0.380 2.360 ;
        RECT  0.100 2.140 1.460 2.300 ;
    END
END AOI12HHD

MACRO AOI12KHD
    CLASS CORE ;
    FOREIGN AOI12KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.520 3.900 2.680 ;
        RECT  3.440 2.400 3.900 2.680 ;
        RECT  3.700 1.720 5.100 1.880 ;
        RECT  4.900 0.520 5.100 2.680 ;
        RECT  4.900 0.520 5.260 0.800 ;
        RECT  4.900 2.400 5.260 2.680 ;
        RECT  3.440 0.520 3.900 0.800 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.100 1.960 ;
        RECT  0.820 1.400 1.100 1.680 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.500 1.560 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.780 ;
        RECT  1.640 1.400 1.900 1.680 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.280 2.120 0.400 ;
        RECT  2.880 -0.280 3.160 0.400 ;
        RECT  4.200 -0.280 4.480 0.620 ;
        RECT  5.540 -0.280 5.820 0.400 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  0.980 -0.280 1.260 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.880 2.800 3.160 3.480 ;
        RECT  4.200 2.580 4.480 3.480 ;
        RECT  5.540 2.800 5.820 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  1.740 2.800 2.020 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.440 0.960 2.640 2.120 ;
        RECT  2.440 1.400 2.760 1.680 ;
        RECT  0.620 2.480 2.280 2.640 ;
        RECT  2.120 0.780 2.280 2.640 ;
        RECT  1.460 0.780 1.740 1.020 ;
        RECT  0.100 0.780 2.280 0.940 ;
        RECT  0.100 0.720 0.380 0.940 ;
        RECT  0.100 2.080 0.380 2.360 ;
        RECT  0.100 2.140 1.460 2.300 ;
    END
END AOI12KHD

MACRO AOI13BHD
    CLASS CORE ;
    FOREIGN AOI13BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 2.120 1.020 2.280 ;
        RECT  0.100 0.740 3.100 0.900 ;
        RECT  2.900 0.740 3.100 2.360 ;
        RECT  0.860 0.740 1.020 2.280 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AOI13BHD

MACRO AOI13EHD
    CLASS CORE ;
    FOREIGN AOI13EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.460 4.700 2.740 ;
        RECT  4.480 2.460 4.700 2.740 ;
        RECT  4.480 0.460 4.700 0.740 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.860 -0.280 4.140 0.400 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.860 2.800 4.140 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 2.060 3.500 2.340 ;
        RECT  3.300 0.860 3.500 2.340 ;
        RECT  3.300 1.400 3.580 1.680 ;
        RECT  3.280 0.860 3.500 1.140 ;
        RECT  0.100 2.120 1.020 2.280 ;
        RECT  0.860 0.740 1.020 2.280 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AOI13EHD

MACRO AOI13HHD
    CLASS CORE ;
    FOREIGN AOI13HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.520 4.700 2.680 ;
        RECT  4.260 2.400 4.700 2.680 ;
        RECT  4.260 0.520 4.700 0.800 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.700 -0.280 3.980 0.400 ;
        RECT  4.820 -0.280 5.100 0.400 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.700 2.800 3.980 3.480 ;
        RECT  4.820 2.800 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.300 1.400 3.580 1.680 ;
        RECT  3.280 0.460 3.500 0.740 ;
        RECT  0.100 2.120 1.020 2.280 ;
        RECT  0.860 0.740 1.020 2.280 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AOI13HHD

MACRO AOI13KHD
    CLASS CORE ;
    FOREIGN AOI13KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.520 4.700 2.680 ;
        RECT  4.260 2.400 4.700 2.680 ;
        RECT  4.500 1.300 5.500 1.500 ;
        RECT  5.300 0.520 5.500 2.680 ;
        RECT  5.300 0.520 5.660 0.800 ;
        RECT  5.300 2.400 5.660 2.680 ;
        RECT  4.260 0.520 4.700 0.800 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.400 2.700 1.960 ;
        RECT  2.380 1.400 2.700 1.680 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.900 1.360 2.060 1.640 ;
        RECT  1.700 1.060 1.900 1.560 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.060 1.500 1.560 ;
        RECT  1.220 1.360 1.380 1.640 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.380 1.340 0.700 1.620 ;
        RECT  0.500 1.100 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.700 -0.280 3.980 0.400 ;
        RECT  4.820 -0.280 5.100 0.400 ;
        RECT  5.940 -0.280 6.220 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.700 -0.280 0.980 0.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 2.800 2.940 3.480 ;
        RECT  3.700 2.800 3.980 3.480 ;
        RECT  4.820 2.800 5.100 3.480 ;
        RECT  5.940 2.800 6.220 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  1.540 2.800 1.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 2.460 3.500 2.740 ;
        RECT  3.300 0.460 3.500 2.740 ;
        RECT  3.300 1.400 3.580 1.680 ;
        RECT  3.280 0.460 3.500 0.740 ;
        RECT  0.100 2.120 1.020 2.280 ;
        RECT  0.860 0.740 1.020 2.280 ;
        RECT  2.920 0.740 3.080 1.720 ;
        RECT  0.100 0.740 3.080 0.900 ;
        RECT  0.980 2.480 2.380 2.640 ;
    END
END AOI13KHD

MACRO AOI2222CHD
    CLASS CORE ;
    FOREIGN AOI2222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.880 0.860 7.100 2.280 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        RECT  3.260 1.340 3.500 1.620 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.370 4.740 1.650 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  6.100 -0.280 6.380 0.400 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.930 2.800 5.210 3.480 ;
        RECT  6.260 2.800 6.540 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.650 2.120 6.700 2.280 ;
        RECT  6.540 0.600 6.700 2.280 ;
        RECT  5.650 1.960 5.930 2.280 ;
        RECT  5.020 0.600 6.700 0.760 ;
        RECT  2.720 2.600 4.740 2.760 ;
        RECT  4.580 2.300 4.740 2.760 ;
        RECT  2.720 2.120 2.880 2.760 ;
        RECT  4.580 2.300 5.490 2.460 ;
        RECT  5.330 1.640 5.490 2.460 ;
        RECT  1.100 2.120 2.880 2.280 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.330 1.640 6.010 1.800 ;
        RECT  5.730 1.520 6.010 1.800 ;
        RECT  0.580 0.920 1.880 1.080 ;
        RECT  3.540 1.960 5.160 2.120 ;
        RECT  5.000 0.920 5.160 2.120 ;
        RECT  5.000 1.200 5.410 1.460 ;
        RECT  3.020 0.920 5.160 1.080 ;
        RECT  2.540 0.600 4.820 0.760 ;
        RECT  3.060 2.280 4.420 2.440 ;
        RECT  3.060 2.220 3.340 2.440 ;
        RECT  0.100 0.600 2.340 0.760 ;
        RECT  0.620 2.440 1.940 2.600 ;
    END
END AOI2222CHD

MACRO AOI2222EHD
    CLASS CORE ;
    FOREIGN AOI2222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.880 0.920 7.100 2.280 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        RECT  3.260 1.340 3.500 1.620 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.370 4.740 1.650 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  6.100 -0.280 6.380 0.400 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.890 2.800 5.170 3.480 ;
        RECT  6.260 2.800 6.540 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.650 2.320 6.700 2.480 ;
        RECT  6.540 0.600 6.700 2.480 ;
        RECT  5.650 2.160 5.930 2.480 ;
        RECT  5.020 0.600 6.700 0.760 ;
        RECT  2.720 2.280 5.490 2.440 ;
        RECT  5.330 1.830 5.490 2.440 ;
        RECT  1.100 2.120 2.880 2.280 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.330 1.830 5.950 1.990 ;
        RECT  5.790 1.460 5.950 1.990 ;
        RECT  0.580 0.920 1.880 1.080 ;
        RECT  3.540 1.960 5.160 2.120 ;
        RECT  5.000 0.920 5.160 2.120 ;
        RECT  5.000 1.400 5.410 1.560 ;
        RECT  3.020 0.920 5.160 1.080 ;
        RECT  2.540 0.600 4.820 0.760 ;
        RECT  3.020 2.600 4.420 2.760 ;
        RECT  0.100 0.600 2.340 0.760 ;
        RECT  0.620 2.440 1.940 2.600 ;
    END
END AOI2222EHD

MACRO AOI2222HHD
    CLASS CORE ;
    FOREIGN AOI2222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.900 7.500 2.300 ;
        RECT  6.700 2.100 7.500 2.300 ;
        RECT  6.700 0.900 7.500 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        RECT  3.260 1.340 3.500 1.620 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.370 4.740 1.650 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  6.040 -0.280 6.320 0.400 ;
        RECT  7.220 -0.280 7.500 0.580 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.940 2.800 5.220 3.480 ;
        RECT  6.140 2.800 6.420 3.480 ;
        RECT  7.220 2.620 7.500 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.580 2.240 6.540 2.400 ;
        RECT  6.380 0.600 6.540 2.400 ;
        RECT  5.580 2.160 5.860 2.400 ;
        RECT  5.020 0.600 6.540 0.760 ;
        RECT  2.720 2.280 5.420 2.440 ;
        RECT  5.260 1.830 5.420 2.440 ;
        RECT  1.100 2.120 2.880 2.280 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.260 1.830 5.950 1.990 ;
        RECT  5.790 1.460 5.950 1.990 ;
        RECT  0.580 0.920 1.880 1.080 ;
        RECT  3.540 1.960 5.100 2.120 ;
        RECT  4.940 0.920 5.100 2.120 ;
        RECT  4.940 1.400 5.410 1.560 ;
        RECT  3.020 0.920 5.100 1.080 ;
        RECT  2.540 0.600 4.820 0.760 ;
        RECT  3.020 2.600 4.420 2.760 ;
        RECT  0.100 0.600 2.340 0.760 ;
        RECT  0.620 2.440 1.940 2.600 ;
    END
END AOI2222HHD

MACRO AOI2222KHD
    CLASS CORE ;
    FOREIGN AOI2222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.900 9.900 2.300 ;
        RECT  8.060 2.100 9.900 2.300 ;
        RECT  8.060 0.900 9.900 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.760 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.370 4.740 1.650 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        RECT  2.780 1.390 3.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.940 -0.280 4.220 0.400 ;
        RECT  5.020 -0.280 5.300 0.760 ;
        RECT  7.500 -0.280 7.780 0.400 ;
        RECT  8.580 -0.280 8.860 0.580 ;
        RECT  9.620 -0.280 9.900 0.580 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 2.440 2.520 3.480 ;
        RECT  4.640 2.740 4.800 3.480 ;
        RECT  5.960 2.800 6.240 3.480 ;
        RECT  7.500 2.800 7.780 3.480 ;
        RECT  8.580 2.620 8.860 3.480 ;
        RECT  9.620 2.620 9.900 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.360 2.160 7.900 2.320 ;
        RECT  7.740 0.600 7.900 2.320 ;
        RECT  5.900 0.600 7.900 0.760 ;
        RECT  1.100 2.120 2.780 2.280 ;
        RECT  5.000 1.340 5.160 2.120 ;
        RECT  2.620 1.960 5.160 2.120 ;
        RECT  1.720 0.920 1.880 2.280 ;
        RECT  5.000 1.780 6.880 1.940 ;
        RECT  6.720 1.340 6.880 1.940 ;
        RECT  5.000 1.340 5.240 1.620 ;
        RECT  0.580 0.920 1.880 1.080 ;
        RECT  6.400 2.480 6.680 2.760 ;
        RECT  5.000 2.480 6.680 2.640 ;
        RECT  5.000 2.280 5.160 2.640 ;
        RECT  3.440 2.280 5.160 2.440 ;
        RECT  6.220 0.920 6.380 1.620 ;
        RECT  3.020 0.920 6.380 1.080 ;
        RECT  2.540 0.600 4.820 0.760 ;
        RECT  2.920 2.600 4.320 2.760 ;
        RECT  0.100 0.600 2.340 0.760 ;
        RECT  0.620 2.440 1.940 2.600 ;
    END
END AOI2222KHD

MACRO AOI222BHD
    CLASS CORE ;
    FOREIGN AOI222BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.820 4.300 2.320 ;
        RECT  3.500 2.120 4.300 2.320 ;
        RECT  0.100 0.820 4.300 0.980 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.370 2.820 1.650 ;
        RECT  2.500 1.250 2.700 1.890 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.250 2.300 1.890 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.250 3.500 1.890 ;
        RECT  3.220 1.370 3.500 1.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.250 3.900 1.890 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 -0.280 3.260 0.660 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  1.080 -0.280 1.720 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.290 2.440 1.570 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.940 2.600 4.300 2.760 ;
        RECT  1.940 2.450 2.220 2.760 ;
        RECT  0.580 2.120 2.780 2.280 ;
    END
END AOI222BHD

MACRO AOI222EHD
    CLASS CORE ;
    FOREIGN AOI222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.680 0.520 5.900 2.680 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.240 3.900 1.880 ;
        RECT  3.640 1.370 3.900 1.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.860 -0.280 4.140 0.400 ;
        RECT  5.160 -0.280 5.320 0.640 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.220 2.800 2.940 3.480 ;
        RECT  3.880 2.800 4.160 3.480 ;
        RECT  5.060 2.800 5.340 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.100 2.600 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.460 2.220 5.500 2.380 ;
        RECT  5.340 1.020 5.500 2.380 ;
        RECT  4.760 1.020 5.500 1.180 ;
        RECT  3.200 2.320 4.280 2.480 ;
        RECT  4.120 1.880 4.280 2.480 ;
        RECT  4.120 1.880 4.600 2.040 ;
        RECT  4.440 0.600 4.600 2.040 ;
        RECT  4.440 1.430 4.860 1.590 ;
        RECT  2.730 0.600 4.600 0.760 ;
        RECT  1.100 2.280 2.680 2.440 ;
        RECT  2.520 0.920 2.680 2.440 ;
        RECT  4.120 0.920 4.280 1.660 ;
        RECT  0.580 0.920 4.280 1.080 ;
        RECT  0.100 0.600 2.500 0.760 ;
        RECT  0.620 2.600 1.980 2.760 ;
        RECT  0.620 2.540 0.900 2.760 ;
    END
END AOI222EHD

MACRO AOI222HHD
    CLASS CORE ;
    FOREIGN AOI222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.900 6.300 2.300 ;
        RECT  5.500 2.100 6.300 2.300 ;
        RECT  5.500 0.900 6.300 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.370 3.680 1.650 ;
        RECT  3.300 1.240 3.500 1.880 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.760 -0.280 4.040 0.400 ;
        RECT  5.040 -0.280 5.200 0.640 ;
        RECT  6.020 -0.280 6.300 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.220 2.800 2.860 3.480 ;
        RECT  3.760 2.800 4.040 3.480 ;
        RECT  4.940 2.800 5.220 3.480 ;
        RECT  6.020 2.620 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.100 2.600 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.340 2.480 5.300 2.640 ;
        RECT  5.140 1.020 5.300 2.640 ;
        RECT  4.640 1.020 5.300 1.180 ;
        RECT  3.160 2.160 4.480 2.320 ;
        RECT  4.320 0.600 4.480 2.320 ;
        RECT  4.320 1.430 4.740 1.590 ;
        RECT  2.730 0.600 4.480 0.760 ;
        RECT  1.100 2.280 2.680 2.440 ;
        RECT  2.520 0.920 2.680 2.440 ;
        RECT  4.000 0.920 4.160 1.690 ;
        RECT  0.580 0.920 4.160 1.080 ;
        RECT  0.100 0.600 2.500 0.760 ;
        RECT  0.580 2.600 1.980 2.760 ;
    END
END AOI222HHD

MACRO AOI222KHD
    CLASS CORE ;
    FOREIGN AOI222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.900 8.700 2.300 ;
        RECT  6.860 2.100 8.700 2.300 ;
        RECT  6.860 0.900 8.700 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.370 3.680 1.650 ;
        RECT  3.300 1.240 3.500 1.880 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.880 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.760 -0.280 4.040 0.400 ;
        RECT  5.700 -0.280 5.980 0.400 ;
        RECT  7.380 -0.280 7.660 0.580 ;
        RECT  8.420 -0.280 8.700 0.580 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 2.800 2.650 3.480 ;
        RECT  3.660 2.800 3.940 3.480 ;
        RECT  4.780 2.800 5.060 3.480 ;
        RECT  6.340 2.620 6.620 3.480 ;
        RECT  7.380 2.620 7.660 3.480 ;
        RECT  8.420 2.620 8.700 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.600 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.180 2.100 6.700 2.260 ;
        RECT  6.540 0.620 6.700 2.260 ;
        RECT  4.640 0.620 6.700 0.780 ;
        RECT  1.100 2.120 2.680 2.280 ;
        RECT  2.520 0.920 2.680 2.280 ;
        RECT  4.000 1.780 5.700 1.940 ;
        RECT  5.540 1.340 5.700 1.940 ;
        RECT  4.000 0.920 4.160 1.940 ;
        RECT  0.580 0.920 4.160 1.080 ;
        RECT  5.220 2.480 5.500 2.760 ;
        RECT  3.720 2.480 5.500 2.640 ;
        RECT  3.100 2.380 3.880 2.540 ;
        RECT  4.960 1.010 5.120 1.620 ;
        RECT  4.320 1.010 5.120 1.170 ;
        RECT  4.320 0.600 4.480 1.170 ;
        RECT  2.700 0.600 4.480 0.760 ;
        RECT  0.100 0.600 2.500 0.760 ;
        RECT  0.620 2.600 1.980 2.760 ;
        RECT  0.620 2.540 0.900 2.760 ;
    END
END AOI222KHD

MACRO AOI22BHD
    CLASS CORE ;
    FOREIGN AOI22BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.920 2.700 2.280 ;
        RECT  1.100 2.120 2.700 2.280 ;
        RECT  0.580 0.920 2.700 1.080 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.340 1.650 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  1.560 -0.280 1.840 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 2.440 2.620 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 0.600 2.620 0.760 ;
        RECT  0.620 2.440 1.940 2.600 ;
    END
END AOI22BHD

MACRO AOI22EHD
    CLASS CORE ;
    FOREIGN AOI22EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 0.520 4.300 2.680 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.520 -0.280 3.680 0.820 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  1.560 -0.280 1.840 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.620 2.480 3.480 ;
        RECT  3.520 2.380 3.680 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.860 1.900 3.020 2.540 ;
        RECT  2.860 1.900 3.900 2.060 ;
        RECT  3.740 1.020 3.900 2.060 ;
        RECT  2.800 1.020 3.900 1.180 ;
        RECT  1.100 2.280 2.640 2.440 ;
        RECT  2.480 0.880 2.640 2.440 ;
        RECT  2.480 1.430 3.260 1.590 ;
        RECT  0.580 0.880 2.640 1.040 ;
        RECT  0.100 0.560 2.600 0.720 ;
        RECT  0.620 2.600 1.940 2.760 ;
        RECT  0.620 2.540 0.900 2.760 ;
    END
END AOI22EHD

MACRO AOI22HHD
    CLASS CORE ;
    FOREIGN AOI22HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.900 4.700 2.300 ;
        RECT  3.900 2.100 4.700 2.300 ;
        RECT  3.900 0.900 4.700 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.380 -0.280 3.660 0.580 ;
        RECT  4.420 -0.280 4.700 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  1.560 -0.280 1.840 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.420 2.480 3.480 ;
        RECT  3.440 2.380 3.600 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.920 1.900 3.080 2.540 ;
        RECT  2.920 1.900 3.740 2.060 ;
        RECT  3.580 1.020 3.740 2.060 ;
        RECT  2.860 1.020 3.740 1.180 ;
        RECT  1.100 2.100 2.700 2.260 ;
        RECT  2.540 0.920 2.700 2.260 ;
        RECT  2.540 1.430 3.320 1.590 ;
        RECT  0.580 0.920 2.700 1.080 ;
        RECT  0.100 0.600 2.600 0.760 ;
        RECT  0.620 2.420 1.980 2.580 ;
    END
END AOI22HHD

MACRO AOI22KHD
    CLASS CORE ;
    FOREIGN AOI22KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.860 5.900 2.300 ;
        RECT  4.050 2.100 5.900 2.300 ;
        RECT  4.050 0.860 5.900 1.060 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.880 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.880 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.530 -0.280 3.810 0.580 ;
        RECT  4.580 -0.280 4.860 0.580 ;
        RECT  5.620 -0.280 5.900 0.580 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  1.560 -0.280 1.840 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 2.420 2.600 3.480 ;
        RECT  3.530 2.620 3.810 3.480 ;
        RECT  4.580 2.620 4.860 3.480 ;
        RECT  5.620 2.620 5.900 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.070 1.900 3.230 2.540 ;
        RECT  3.070 1.900 3.890 2.060 ;
        RECT  3.730 1.020 3.890 2.060 ;
        RECT  3.010 1.020 3.890 1.180 ;
        RECT  1.100 2.100 2.700 2.260 ;
        RECT  2.540 0.920 2.700 2.260 ;
        RECT  2.540 1.430 3.470 1.590 ;
        RECT  0.580 0.920 2.700 1.080 ;
        RECT  0.100 0.600 2.600 0.760 ;
        RECT  0.100 0.560 0.380 0.760 ;
        RECT  0.580 2.420 1.980 2.580 ;
    END
END AOI22KHD

MACRO BHD1HD
    CLASS CORE ;
    FOREIGN BHD1HD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN H
        DIRECTION INOUT ;
        PORT
        LAYER metal1 ;
        RECT  0.800 1.240 1.000 2.450 ;
        RECT  2.780 0.960 3.100 1.240 ;
        RECT  2.780 1.840 3.100 2.120 ;
        RECT  2.900 0.920 3.100 2.450 ;
        RECT  0.800 2.290 3.100 2.450 ;
        RECT  0.720 1.370 1.000 1.650 ;
        END
    END H
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.620 -0.280 2.060 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.620 2.620 2.060 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 0.880 0.320 2.160 ;
        RECT  2.220 0.880 2.380 1.660 ;
        RECT  0.160 0.880 2.380 1.040 ;
    END
END BHD1HD

MACRO BUFBEHD
    CLASS CORE ;
    FOREIGN BUFBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.760 1.900 2.360 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.920 2.300 1.960 ;
        RECT  2.100 0.920 3.080 1.080 ;
        RECT  2.920 0.920 3.080 1.740 ;
        RECT  2.920 1.460 3.180 1.740 ;
        RECT  2.060 1.460 2.300 1.740 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 -0.280 2.980 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 2.800 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 1.960 3.500 2.240 ;
        RECT  3.340 0.560 3.500 2.240 ;
        RECT  1.380 0.440 1.540 1.510 ;
        RECT  3.280 0.960 3.500 1.240 ;
        RECT  2.120 0.560 3.500 0.720 ;
        RECT  1.380 0.440 2.280 0.600 ;
        RECT  1.320 2.520 2.280 2.680 ;
        RECT  2.120 2.120 2.280 2.680 ;
        RECT  1.320 2.120 1.480 2.680 ;
        RECT  2.120 2.120 2.700 2.280 ;
        RECT  2.540 1.460 2.700 2.280 ;
        RECT  0.100 2.120 1.480 2.280 ;
        RECT  0.900 1.370 1.060 2.280 ;
        RECT  0.100 0.840 0.260 2.280 ;
        RECT  0.100 0.840 0.320 1.120 ;
    END
END BUFBEHD

MACRO BUFBHHD
    CLASS CORE ;
    FOREIGN BUFBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.400 2.120 4.300 2.280 ;
        RECT  4.100 0.740 4.300 2.360 ;
        RECT  3.500 0.740 4.300 0.900 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.540 -0.280 1.820 0.400 ;
        RECT  2.900 -0.280 3.180 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.600 -0.280 0.880 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 2.800 2.120 3.480 ;
        RECT  3.040 2.560 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.320 1.900 1.700 2.060 ;
        RECT  1.320 0.560 1.480 2.060 ;
        RECT  3.180 1.200 3.940 1.360 ;
        RECT  3.180 0.560 3.340 1.360 ;
        RECT  1.160 0.740 1.480 1.020 ;
        RECT  1.320 0.560 3.340 0.720 ;
        RECT  2.480 0.920 2.640 2.120 ;
        RECT  2.480 1.520 3.540 1.680 ;
        RECT  1.980 0.920 2.640 1.080 ;
        RECT  2.600 2.480 2.880 2.690 ;
        RECT  1.320 2.480 2.880 2.640 ;
        RECT  1.320 2.300 1.480 2.640 ;
        RECT  0.100 2.300 1.480 2.460 ;
        RECT  0.100 1.840 0.320 2.460 ;
        RECT  0.100 0.910 0.260 2.460 ;
        RECT  0.100 0.910 0.320 1.190 ;
    END
END BUFBHHD

MACRO BUFBIHD
    CLASS CORE ;
    FOREIGN BUFBIHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.500 0.740 4.820 0.900 ;
        RECT  3.500 2.120 4.980 2.280 ;
        RECT  4.500 0.740 4.700 2.360 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.540 -0.280 1.820 0.400 ;
        RECT  2.900 -0.280 3.180 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.600 -0.280 0.880 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 2.800 2.120 3.480 ;
        RECT  3.040 2.560 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.320 1.900 1.700 2.060 ;
        RECT  1.320 0.560 1.480 2.060 ;
        RECT  3.180 1.250 4.080 1.410 ;
        RECT  3.180 0.560 3.340 1.410 ;
        RECT  1.160 0.740 1.480 1.020 ;
        RECT  1.320 0.560 3.340 0.720 ;
        RECT  2.480 0.920 2.640 2.120 ;
        RECT  2.480 1.690 3.600 1.850 ;
        RECT  1.960 0.920 2.640 1.080 ;
        RECT  2.600 2.480 2.880 2.690 ;
        RECT  1.320 2.480 2.880 2.640 ;
        RECT  1.320 2.300 1.480 2.640 ;
        RECT  0.100 2.300 1.480 2.460 ;
        RECT  0.100 1.840 0.320 2.460 ;
        RECT  0.100 0.910 0.260 2.460 ;
        RECT  0.100 0.910 0.320 1.190 ;
    END
END BUFBIHD

MACRO BUFBKHD
    CLASS CORE ;
    FOREIGN BUFBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.500 0.740 4.980 0.900 ;
        RECT  3.410 2.120 5.090 2.280 ;
        RECT  4.500 0.740 4.700 2.360 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END EB
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.540 -0.280 1.820 0.400 ;
        RECT  2.900 -0.280 3.180 0.400 ;
        RECT  4.100 -0.280 4.380 0.400 ;
        RECT  5.220 -0.280 5.500 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.600 -0.280 0.880 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 2.800 2.120 3.480 ;
        RECT  3.040 2.560 3.260 3.480 ;
        RECT  4.100 2.800 4.380 3.480 ;
        RECT  5.220 2.620 5.500 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.320 1.900 1.700 2.060 ;
        RECT  1.320 0.560 1.480 2.060 ;
        RECT  2.920 1.200 3.840 1.360 ;
        RECT  2.920 0.560 3.080 1.360 ;
        RECT  1.160 0.740 1.480 1.020 ;
        RECT  1.320 0.560 3.080 0.720 ;
        RECT  2.480 0.920 2.640 2.120 ;
        RECT  2.480 1.520 3.420 1.680 ;
        RECT  1.970 0.920 2.640 1.080 ;
        RECT  2.600 2.480 2.880 2.690 ;
        RECT  1.320 2.480 2.880 2.640 ;
        RECT  1.320 2.300 1.480 2.640 ;
        RECT  0.100 2.300 1.480 2.460 ;
        RECT  0.100 1.840 0.320 2.460 ;
        RECT  0.100 0.910 0.260 2.460 ;
        RECT  0.100 0.910 0.320 1.190 ;
    END
END BUFBKHD

MACRO BUFCHD
    CLASS CORE ;
    FOREIGN BUFCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.660 1.500 2.440 ;
        RECT  1.280 2.160 1.500 2.440 ;
        RECT  1.280 0.660 1.500 0.940 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.210 0.380 2.430 ;
        RECT  0.100 2.210 1.080 2.370 ;
        RECT  0.920 0.720 1.080 2.370 ;
        RECT  0.920 1.460 1.140 1.740 ;
        RECT  0.100 0.720 1.080 0.880 ;
        RECT  0.100 0.660 0.380 0.880 ;
    END
END BUFCHD

MACRO BUFCKEHD
    CLASS CORE ;
    FOREIGN BUFCKEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 0.580 1.480 2.740 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.230 1.080 2.390 ;
        RECT  0.920 0.820 1.080 2.390 ;
        RECT  0.100 0.820 1.080 0.980 ;
    END
END BUFCKEHD

MACRO BUFCKGHD
    CLASS CORE ;
    FOREIGN BUFCKGHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.900 2.700 2.300 ;
        RECT  1.900 2.100 2.700 2.300 ;
        RECT  1.860 0.900 2.700 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  1.260 -0.280 1.540 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.280 2.670 1.560 3.480 ;
        RECT  2.420 2.530 2.700 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 2.330 1.540 2.490 ;
        RECT  1.380 0.820 1.540 2.490 ;
        RECT  0.620 0.820 1.540 0.980 ;
    END
END BUFCKGHD

MACRO BUFCKHHD
    CLASS CORE ;
    FOREIGN BUFCKHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.900 2.700 2.300 ;
        RECT  1.900 2.100 2.700 2.300 ;
        RECT  1.820 0.900 2.700 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.370 0.780 1.650 ;
        RECT  0.500 1.320 0.700 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  1.260 -0.280 1.540 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.340 2.800 1.620 3.480 ;
        RECT  2.420 2.620 2.700 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.180 2.560 0.460 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.740 2.370 1.600 2.530 ;
        RECT  1.440 0.850 1.600 2.530 ;
        RECT  1.440 1.370 1.660 1.650 ;
        RECT  0.620 0.850 1.600 1.010 ;
    END
END BUFCKHHD

MACRO BUFCKIHD
    CLASS CORE ;
    FOREIGN BUFCKIHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.840 1.960 2.030 2.240 ;
        RECT  1.870 0.860 2.080 1.140 ;
        RECT  2.880 0.830 3.080 1.110 ;
        RECT  1.870 1.420 3.080 1.680 ;
        RECT  2.920 0.830 3.080 2.350 ;
        RECT  2.880 2.070 3.080 2.350 ;
        RECT  1.870 0.860 2.030 2.240 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.260 -0.280 2.540 0.400 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  1.260 -0.280 1.540 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.580 1.460 3.480 ;
        RECT  2.300 2.620 2.580 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.100 2.520 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.580 2.260 1.540 2.420 ;
        RECT  1.380 0.850 1.540 2.420 ;
        RECT  0.620 0.850 1.540 1.010 ;
    END
END BUFCKIHD

MACRO BUFCKJHD
    CLASS CORE ;
    FOREIGN BUFCKJHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.240 2.060 2.480 2.340 ;
        RECT  3.280 0.870 3.480 1.150 ;
        RECT  2.320 1.440 3.480 1.740 ;
        RECT  3.320 0.870 3.480 2.340 ;
        RECT  3.280 2.060 3.480 2.340 ;
        RECT  2.320 0.870 2.480 2.340 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.640 ;
        RECT  2.660 -0.280 2.940 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.140 -0.280 0.780 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.520 2.580 1.800 3.480 ;
        RECT  2.700 2.620 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.300 1.360 2.460 ;
        RECT  1.200 0.790 1.360 2.460 ;
        RECT  1.200 1.430 2.120 1.590 ;
    END
END BUFCKJHD

MACRO BUFCKKHD
    CLASS CORE ;
    FOREIGN BUFCKKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 0.860 3.440 2.340 ;
        RECT  3.280 2.060 3.480 2.340 ;
        RECT  4.320 0.860 4.680 1.770 ;
        RECT  3.280 1.370 4.680 1.770 ;
        RECT  4.360 0.860 4.680 2.340 ;
        RECT  3.200 0.860 3.440 1.140 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.320 1.100 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 -0.280 1.740 0.400 ;
        RECT  2.580 -0.280 2.860 0.400 ;
        RECT  3.700 -0.280 3.980 0.640 ;
        RECT  4.820 -0.280 5.100 0.400 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.140 -0.280 0.420 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.480 2.620 1.760 3.480 ;
        RECT  2.740 2.580 3.020 3.480 ;
        RECT  3.780 2.620 4.060 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.180 2.420 0.460 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.920 2.180 2.920 2.340 ;
        RECT  2.760 0.920 2.920 2.340 ;
        RECT  2.760 1.370 3.080 1.650 ;
        RECT  0.860 0.920 2.920 1.080 ;
    END
END BUFCKKHD

MACRO BUFCKLHD
    CLASS CORE ;
    FOREIGN BUFCKLHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.860 0.920 3.020 2.280 ;
        RECT  2.740 2.120 3.020 2.280 ;
        RECT  3.760 0.780 3.920 1.870 ;
        RECT  3.780 1.310 3.940 2.280 ;
        RECT  3.780 2.120 4.060 2.280 ;
        RECT  4.880 0.780 5.040 2.340 ;
        RECT  2.860 1.310 5.080 1.870 ;
        RECT  2.580 0.920 3.020 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.380 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.980 -0.280 2.260 0.400 ;
        RECT  3.140 -0.280 3.420 0.640 ;
        RECT  4.260 -0.280 4.540 0.660 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.860 -0.280 1.140 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.380 1.460 3.480 ;
        RECT  2.220 2.380 2.500 3.480 ;
        RECT  3.260 2.580 3.540 3.480 ;
        RECT  4.300 2.580 4.580 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.380 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 2.020 2.280 2.180 ;
        RECT  2.120 0.600 2.280 2.180 ;
        RECT  2.120 1.430 2.680 1.590 ;
        RECT  0.260 0.600 2.280 0.760 ;
    END
END BUFCKLHD

MACRO BUFCKMHD
    CLASS CORE ;
    FOREIGN BUFCKMHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.420 0.920 3.700 2.340 ;
        RECT  4.340 0.920 4.740 1.080 ;
        RECT  4.460 0.920 4.740 2.340 ;
        RECT  3.420 1.320 5.740 1.880 ;
        RECT  5.460 0.920 5.740 2.340 ;
        RECT  5.460 2.120 5.780 2.280 ;
        RECT  3.220 0.920 3.700 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.430 1.980 1.590 ;
        RECT  1.300 1.320 1.500 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.450 -0.280 1.730 0.400 ;
        RECT  2.620 -0.280 2.900 0.400 ;
        RECT  3.780 -0.280 4.060 0.640 ;
        RECT  4.900 -0.280 5.180 0.660 ;
        RECT  6.020 -0.280 6.300 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.620 2.140 3.480 ;
        RECT  2.900 2.620 3.180 3.480 ;
        RECT  3.940 2.620 4.220 3.480 ;
        RECT  4.980 2.620 5.260 3.480 ;
        RECT  6.020 2.620 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.820 2.620 1.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.260 2.300 2.600 2.460 ;
        RECT  2.440 2.020 2.600 2.460 ;
        RECT  0.260 2.240 0.540 2.460 ;
        RECT  2.440 2.020 3.040 2.180 ;
        RECT  2.880 0.600 3.040 2.180 ;
        RECT  2.760 1.430 3.040 1.590 ;
        RECT  0.860 0.600 3.040 0.760 ;
    END
END BUFCKMHD

MACRO BUFCKNHD
    CLASS CORE ;
    FOREIGN BUFCKNHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.740 0.920 5.020 2.340 ;
        RECT  5.580 0.920 6.060 1.080 ;
        RECT  5.780 0.920 6.060 2.340 ;
        RECT  6.700 0.920 7.100 1.080 ;
        RECT  6.820 0.920 7.100 2.340 ;
        RECT  7.820 0.920 8.140 1.080 ;
        RECT  4.740 1.350 8.140 1.910 ;
        RECT  7.860 0.920 8.140 2.340 ;
        RECT  4.460 0.920 5.020 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.430 2.390 1.590 ;
        RECT  1.700 1.320 1.900 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.760 -0.280 3.040 0.400 ;
        RECT  3.900 -0.280 4.180 0.400 ;
        RECT  5.020 -0.280 5.300 0.640 ;
        RECT  6.140 -0.280 6.420 0.660 ;
        RECT  7.260 -0.280 7.540 0.660 ;
        RECT  8.420 -0.280 8.700 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  1.610 -0.280 1.890 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.940 2.620 2.220 3.480 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.220 2.580 4.500 3.480 ;
        RECT  5.260 2.620 5.540 3.480 ;
        RECT  6.300 2.620 6.580 3.480 ;
        RECT  7.340 2.620 7.620 3.480 ;
        RECT  8.420 2.620 8.700 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.900 2.620 1.180 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.280 2.300 3.720 2.460 ;
        RECT  3.560 0.630 3.720 2.460 ;
        RECT  3.560 1.430 4.280 1.590 ;
        RECT  0.900 0.630 3.720 0.790 ;
    END
END BUFCKNHD

MACRO BUFCKQHD
    CLASS CORE ;
    FOREIGN BUFCKQHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.470 0.920 14.710 2.110 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.660 1.430 3.550 1.590 ;
        RECT  1.700 1.320 1.900 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 -0.280 3.260 0.400 ;
        RECT  4.140 -0.280 4.420 0.400 ;
        RECT  4.910 -0.280 5.190 0.400 ;
        RECT  6.030 -0.280 6.310 0.400 ;
        RECT  7.150 -0.280 7.430 0.400 ;
        RECT  8.270 -0.280 8.550 0.400 ;
        RECT  9.390 -0.280 9.670 0.400 ;
        RECT  10.510 -0.280 10.790 0.400 ;
        RECT  11.630 -0.280 11.910 0.400 ;
        RECT  12.750 -0.280 13.030 0.400 ;
        RECT  13.870 -0.280 14.150 0.400 ;
        RECT  14.990 -0.280 15.270 0.400 ;
        RECT  0.000 -0.280 15.600 0.280 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.820 2.620 2.100 3.480 ;
        RECT  2.860 2.620 3.140 3.480 ;
        RECT  3.900 2.620 4.180 3.480 ;
        RECT  5.230 2.580 5.510 3.480 ;
        RECT  6.270 2.620 6.550 3.480 ;
        RECT  7.310 2.620 7.590 3.480 ;
        RECT  8.350 2.620 8.630 3.480 ;
        RECT  9.390 2.620 9.670 3.480 ;
        RECT  10.430 2.620 10.710 3.480 ;
        RECT  11.470 2.620 11.750 3.480 ;
        RECT  12.510 2.620 12.790 3.480 ;
        RECT  13.550 2.620 13.830 3.480 ;
        RECT  14.590 2.580 14.870 3.480 ;
        RECT  0.000 2.920 15.600 3.480 ;
        RECT  0.780 2.620 1.060 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.220 2.220 4.850 2.460 ;
        RECT  4.610 0.660 4.850 2.460 ;
        RECT  4.610 1.390 5.250 1.630 ;
        RECT  1.300 0.660 4.850 0.900 ;
    END
END BUFCKQHD

MACRO BUFDHD
    CLASS CORE ;
    FOREIGN BUFDHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.660 1.500 2.440 ;
        RECT  1.280 2.160 1.500 2.440 ;
        RECT  1.280 0.660 1.500 0.940 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.210 0.380 2.430 ;
        RECT  0.100 2.210 1.080 2.370 ;
        RECT  0.920 0.720 1.080 2.370 ;
        RECT  0.920 1.460 1.140 1.740 ;
        RECT  0.100 0.720 1.080 0.880 ;
        RECT  0.100 0.660 0.380 0.880 ;
    END
END BUFDHD

MACRO BUFEHD
    CLASS CORE ;
    FOREIGN BUFEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.660 1.500 2.440 ;
        RECT  1.280 2.160 1.500 2.440 ;
        RECT  1.280 0.660 1.500 0.940 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.210 0.380 2.430 ;
        RECT  0.100 2.210 1.080 2.370 ;
        RECT  0.920 0.720 1.080 2.370 ;
        RECT  0.920 1.460 1.140 1.740 ;
        RECT  0.100 0.720 1.080 0.880 ;
        RECT  0.100 0.660 0.380 0.880 ;
    END
END BUFEHD

MACRO BUFGHD
    CLASS CORE ;
    FOREIGN BUFGHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.660 1.500 2.440 ;
        RECT  1.160 2.160 1.500 2.440 ;
        RECT  1.160 0.660 1.500 0.940 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.680 -0.280 1.840 0.910 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.680 2.250 1.840 3.480 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.120 0.380 2.340 ;
        RECT  0.100 2.120 0.980 2.280 ;
        RECT  0.820 0.860 0.980 2.280 ;
        RECT  0.100 0.860 0.980 1.080 ;
    END
END BUFGHD

MACRO BUFHHD
    CLASS CORE ;
    FOREIGN BUFHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.660 1.500 2.440 ;
        RECT  1.160 2.160 1.500 2.440 ;
        RECT  1.160 0.660 1.500 0.940 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.680 -0.280 1.840 0.770 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.680 2.360 1.840 3.480 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.120 0.380 2.340 ;
        RECT  0.100 2.120 0.980 2.280 ;
        RECT  0.820 0.860 0.980 2.280 ;
        RECT  0.100 0.860 0.980 1.080 ;
    END
END BUFHHD

MACRO BUFIHD
    CLASS CORE ;
    FOREIGN BUFIHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 2.120 1.520 2.340 ;
        RECT  1.240 0.920 2.700 1.080 ;
        RECT  1.240 2.120 2.700 2.280 ;
        RECT  2.480 0.840 2.700 1.120 ;
        RECT  2.480 2.060 2.700 2.340 ;
        RECT  2.500 0.840 2.700 2.360 ;
        RECT  1.240 0.860 1.520 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.760 -0.280 2.040 0.580 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.760 2.620 2.040 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.120 0.380 2.340 ;
        RECT  0.100 2.120 1.080 2.280 ;
        RECT  0.920 0.860 1.080 2.280 ;
        RECT  0.100 0.860 1.080 1.080 ;
    END
END BUFIHD

MACRO BUFJHD
    CLASS CORE ;
    FOREIGN BUFJHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 2.120 2.700 2.280 ;
        RECT  2.480 0.840 2.700 1.120 ;
        RECT  2.480 2.060 2.700 2.340 ;
        RECT  2.500 0.840 2.700 2.360 ;
        RECT  1.280 0.920 2.700 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.580 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.720 -0.280 1.000 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.620 2.140 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.720 2.620 1.000 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.120 0.380 2.340 ;
        RECT  0.100 2.120 1.080 2.280 ;
        RECT  0.920 0.860 1.080 2.280 ;
        RECT  0.100 0.860 1.080 1.080 ;
    END
END BUFJHD

MACRO BUFKHD
    CLASS CORE ;
    FOREIGN BUFKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 2.120 1.940 2.340 ;
        RECT  1.660 0.920 3.100 1.080 ;
        RECT  1.660 2.120 3.100 2.280 ;
        RECT  2.900 0.840 3.100 2.360 ;
        RECT  1.660 0.860 1.940 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  2.180 -0.280 2.460 0.580 ;
        RECT  3.220 -0.280 3.500 0.580 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.100 -0.280 0.380 1.080 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.620 1.420 3.480 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  3.220 2.620 3.500 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.180 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.580 2.120 1.500 2.280 ;
        RECT  1.340 0.920 1.500 2.280 ;
        RECT  0.580 0.920 1.500 1.080 ;
    END
END BUFKHD

MACRO BUFLHD
    CLASS CORE ;
    FOREIGN BUFLHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 2.120 1.940 2.340 ;
        RECT  1.660 0.920 3.960 1.080 ;
        RECT  1.660 2.120 3.960 2.280 ;
        RECT  3.700 0.840 3.900 2.360 ;
        RECT  3.700 0.860 3.960 1.140 ;
        RECT  3.700 2.060 3.960 2.340 ;
        RECT  1.660 0.860 1.940 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  2.180 -0.280 2.460 0.580 ;
        RECT  3.220 -0.280 3.500 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 1.080 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.620 1.420 3.480 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  3.220 2.620 3.500 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.180 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.580 2.120 1.500 2.280 ;
        RECT  1.340 0.920 1.500 2.280 ;
        RECT  0.580 0.920 1.500 1.080 ;
    END
END BUFLHD

MACRO BUFMHD
    CLASS CORE ;
    FOREIGN BUFMHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.220 2.120 2.500 2.340 ;
        RECT  2.220 0.920 4.700 1.080 ;
        RECT  2.220 2.120 4.700 2.280 ;
        RECT  4.500 0.840 4.700 2.360 ;
        RECT  2.220 0.860 2.500 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.420 -0.280 1.700 0.780 ;
        RECT  2.740 -0.280 3.020 0.580 ;
        RECT  3.780 -0.280 4.060 0.580 ;
        RECT  4.820 -0.280 5.100 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.420 2.420 1.700 3.480 ;
        RECT  2.740 2.620 3.020 3.480 ;
        RECT  3.780 2.620 4.060 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.560 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.580 2.100 2.060 2.260 ;
        RECT  1.900 0.940 2.060 2.260 ;
        RECT  0.580 0.940 2.060 1.100 ;
    END
END BUFMHD

MACRO BUFNHD
    CLASS CORE ;
    FOREIGN BUFNHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 2.070 2.660 2.340 ;
        RECT  4.070 0.840 4.330 2.360 ;
        RECT  2.380 0.870 5.900 1.130 ;
        RECT  2.380 2.070 5.900 2.330 ;
        RECT  2.380 0.860 2.660 1.130 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.580 ;
        RECT  2.900 -0.280 3.180 0.580 ;
        RECT  3.940 -0.280 4.220 0.580 ;
        RECT  4.980 -0.280 5.260 0.580 ;
        RECT  6.020 -0.280 6.300 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.780 -0.280 1.060 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.620 2.140 3.480 ;
        RECT  2.900 2.620 3.180 3.480 ;
        RECT  3.940 2.620 4.220 3.480 ;
        RECT  4.980 2.620 5.260 3.480 ;
        RECT  6.020 2.620 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.780 2.800 1.060 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.140 2.120 0.420 2.340 ;
        RECT  0.140 2.120 2.220 2.280 ;
        RECT  2.060 0.940 2.220 2.280 ;
        RECT  0.140 0.940 2.220 1.100 ;
    END
END BUFNHD

MACRO BUFQHD
    CLASS CORE ;
    FOREIGN BUFQHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.950 14.100 2.150 ;
        RECT  4.380 1.780 14.100 2.150 ;
        RECT  4.380 0.950 14.100 1.290 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 1.500 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.780 -0.280 2.060 0.580 ;
        RECT  2.820 -0.280 3.100 0.580 ;
        RECT  3.860 -0.280 4.140 0.580 ;
        RECT  4.900 -0.280 5.180 0.580 ;
        RECT  5.940 -0.280 6.220 0.580 ;
        RECT  6.980 -0.280 7.260 0.580 ;
        RECT  8.020 -0.280 8.300 0.580 ;
        RECT  9.060 -0.280 9.340 0.580 ;
        RECT  10.100 -0.280 10.380 0.580 ;
        RECT  11.140 -0.280 11.420 0.580 ;
        RECT  12.180 -0.280 12.460 0.580 ;
        RECT  13.220 -0.280 13.500 0.580 ;
        RECT  14.300 -0.280 14.580 0.400 ;
        RECT  0.000 -0.280 15.200 0.280 ;
        RECT  0.700 -0.280 0.980 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.780 2.620 2.060 3.480 ;
        RECT  2.820 2.620 3.100 3.480 ;
        RECT  3.860 2.620 4.140 3.480 ;
        RECT  4.900 2.620 5.180 3.480 ;
        RECT  5.940 2.620 6.220 3.480 ;
        RECT  6.980 2.620 7.260 3.480 ;
        RECT  8.020 2.620 8.300 3.480 ;
        RECT  9.060 2.620 9.340 3.480 ;
        RECT  10.100 2.620 10.380 3.480 ;
        RECT  11.140 2.620 11.420 3.480 ;
        RECT  12.180 2.620 12.460 3.480 ;
        RECT  13.220 2.620 13.500 3.480 ;
        RECT  14.300 2.800 14.580 3.480 ;
        RECT  0.000 2.920 15.200 3.480 ;
        RECT  0.700 2.800 0.980 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.140 2.120 0.420 2.340 ;
        RECT  0.140 2.120 4.160 2.280 ;
        RECT  4.000 0.920 4.160 2.280 ;
        RECT  4.000 1.460 5.000 1.620 ;
        RECT  0.140 0.920 4.160 1.080 ;
        RECT  0.140 0.860 0.420 1.080 ;
    END
END BUFQHD

MACRO BUFTEHD
    CLASS CORE ;
    FOREIGN BUFTEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.760 1.900 2.360 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.920 2.300 1.960 ;
        RECT  2.100 0.920 3.080 1.080 ;
        RECT  2.920 0.920 3.080 1.740 ;
        RECT  2.920 1.460 3.180 1.740 ;
        RECT  2.060 1.140 2.300 1.420 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 -0.280 2.980 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 2.800 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.280 1.960 3.500 2.240 ;
        RECT  3.340 0.560 3.500 2.240 ;
        RECT  1.380 0.440 1.540 1.740 ;
        RECT  3.280 0.960 3.500 1.240 ;
        RECT  2.120 0.560 3.500 0.720 ;
        RECT  1.380 0.440 2.280 0.600 ;
        RECT  1.320 2.520 2.280 2.680 ;
        RECT  2.120 2.120 2.280 2.680 ;
        RECT  1.320 2.120 1.480 2.680 ;
        RECT  2.120 2.120 2.700 2.280 ;
        RECT  2.540 1.460 2.700 2.280 ;
        RECT  0.100 2.120 1.480 2.280 ;
        RECT  0.900 1.460 1.060 2.280 ;
        RECT  0.100 0.840 0.260 2.280 ;
        RECT  0.100 0.840 0.320 1.120 ;
    END
END BUFTEHD

MACRO BUFTHHD
    CLASS CORE ;
    FOREIGN BUFTHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.740 4.300 2.460 ;
        RECT  3.500 2.300 4.300 2.460 ;
        RECT  3.500 0.740 4.300 0.900 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.820 -0.280 2.100 0.400 ;
        RECT  2.940 -0.280 3.220 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 2.800 1.940 3.480 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.630 2.800 0.910 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.320 2.300 3.080 2.460 ;
        RECT  2.920 1.980 3.080 2.460 ;
        RECT  1.220 2.060 1.480 2.340 ;
        RECT  2.920 1.980 3.940 2.140 ;
        RECT  3.780 1.460 3.940 2.140 ;
        RECT  1.320 0.890 1.480 2.460 ;
        RECT  1.320 0.890 1.700 1.080 ;
        RECT  2.140 1.920 2.660 2.140 ;
        RECT  2.500 0.880 2.660 2.140 ;
        RECT  2.500 1.640 3.460 1.800 ;
        RECT  3.300 1.140 3.460 1.800 ;
        RECT  2.380 0.880 2.660 1.100 ;
        RECT  0.100 2.150 0.320 2.430 ;
        RECT  0.100 0.560 0.260 2.430 ;
        RECT  2.820 0.560 2.980 1.480 ;
        RECT  0.100 0.560 0.320 1.190 ;
        RECT  0.100 0.560 2.980 0.720 ;
    END
END BUFTHHD

MACRO BUFTIHD
    CLASS CORE ;
    FOREIGN BUFTIHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.500 0.740 4.820 0.900 ;
        RECT  3.500 2.300 4.820 2.460 ;
        RECT  4.500 0.740 4.700 2.460 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.820 -0.280 2.100 0.400 ;
        RECT  2.940 -0.280 3.220 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 2.800 1.940 3.480 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.630 2.800 0.910 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.320 2.300 3.080 2.460 ;
        RECT  2.920 1.980 3.080 2.460 ;
        RECT  1.220 2.060 1.480 2.340 ;
        RECT  2.920 1.980 3.940 2.140 ;
        RECT  3.780 1.630 3.940 2.140 ;
        RECT  1.320 0.880 1.480 2.460 ;
        RECT  1.320 0.880 1.700 1.080 ;
        RECT  2.140 1.920 2.660 2.140 ;
        RECT  2.500 0.880 2.660 2.140 ;
        RECT  2.500 1.640 3.480 1.800 ;
        RECT  3.320 1.190 3.480 1.800 ;
        RECT  2.380 0.880 2.660 1.100 ;
        RECT  0.100 2.150 0.320 2.430 ;
        RECT  0.100 0.560 0.260 2.430 ;
        RECT  2.820 0.560 2.980 1.480 ;
        RECT  0.100 0.560 0.320 1.190 ;
        RECT  0.100 0.560 2.980 0.720 ;
    END
END BUFTIHD

MACRO BUFTJHD
    CLASS CORE ;
    FOREIGN BUFTJHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.500 0.740 4.820 0.900 ;
        RECT  3.500 2.300 4.820 2.460 ;
        RECT  4.500 0.740 4.700 2.460 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.820 -0.280 2.100 0.400 ;
        RECT  2.940 -0.280 3.220 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  5.060 -0.280 5.340 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 2.800 1.940 3.480 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  5.060 2.620 5.340 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.630 2.800 0.910 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.320 2.300 3.080 2.460 ;
        RECT  2.920 1.980 3.080 2.460 ;
        RECT  1.220 2.060 1.480 2.340 ;
        RECT  2.920 1.980 3.940 2.140 ;
        RECT  3.780 1.710 3.940 2.140 ;
        RECT  1.320 0.890 1.480 2.460 ;
        RECT  1.320 0.890 1.700 1.080 ;
        RECT  2.140 1.920 2.660 2.140 ;
        RECT  2.500 0.880 2.660 2.140 ;
        RECT  2.500 1.640 3.480 1.800 ;
        RECT  3.320 1.120 3.480 1.800 ;
        RECT  2.380 0.880 2.660 1.100 ;
        RECT  0.100 2.150 0.320 2.430 ;
        RECT  0.100 0.560 0.260 2.430 ;
        RECT  2.820 0.560 2.980 1.480 ;
        RECT  0.100 0.560 0.320 1.190 ;
        RECT  0.100 0.560 2.980 0.720 ;
    END
END BUFTJHD

MACRO BUFTKHD
    CLASS CORE ;
    FOREIGN BUFTKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.660 0.740 4.980 0.900 ;
        RECT  3.660 2.300 4.980 2.460 ;
        RECT  4.500 0.740 4.700 2.460 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.820 -0.280 2.100 0.400 ;
        RECT  3.100 -0.280 3.380 0.400 ;
        RECT  4.180 -0.280 4.460 0.580 ;
        RECT  5.220 -0.280 5.500 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 2.800 1.940 3.480 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.180 2.620 4.460 3.480 ;
        RECT  5.220 2.620 5.500 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.630 2.800 0.910 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.100 1.980 3.120 2.140 ;
        RECT  2.960 0.720 3.120 2.140 ;
        RECT  3.940 1.140 4.220 1.360 ;
        RECT  2.960 1.140 4.220 1.300 ;
        RECT  2.460 0.720 3.120 0.880 ;
        RECT  1.320 2.300 3.480 2.460 ;
        RECT  3.320 1.460 3.480 2.460 ;
        RECT  1.220 2.060 1.480 2.340 ;
        RECT  1.320 0.920 1.480 2.460 ;
        RECT  3.320 1.460 3.540 1.740 ;
        RECT  1.320 0.920 1.700 1.080 ;
        RECT  0.100 2.150 0.320 2.430 ;
        RECT  0.100 0.560 0.260 2.430 ;
        RECT  2.120 1.200 2.800 1.360 ;
        RECT  2.120 0.560 2.280 1.360 ;
        RECT  0.100 0.560 0.320 1.190 ;
        RECT  0.100 0.560 2.280 0.720 ;
    END
END BUFTKHD

MACRO CKLDHD
    CLASS CORE ;
    FOREIGN CKLDHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.320 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        RECT  0.100 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        RECT  0.100 2.440 0.900 3.480 ;
        END
    END VCC
END CKLDHD

MACRO DBAHRBEHD
    CLASS CORE ;
    FOREIGN DBAHRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.340 2.300 1.620 ;
        RECT  2.100 1.000 2.300 1.620 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.520 7.500 2.670 ;
        RECT  7.270 2.390 7.500 2.670 ;
        RECT  7.270 0.520 7.500 0.800 ;
        END
    END QB
    PIN GB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END GB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.340 2.840 1.620 ;
        RECT  2.500 1.000 2.700 1.620 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.850 6.310 1.130 ;
        RECT  6.100 1.840 6.310 2.120 ;
        RECT  6.100 0.850 6.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.760 ;
        RECT  6.690 -0.280 6.970 0.580 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.490 2.470 2.770 3.480 ;
        RECT  5.220 2.740 5.420 3.480 ;
        RECT  6.650 2.800 6.930 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.670 2.300 7.010 2.460 ;
        RECT  6.850 1.420 7.010 2.460 ;
        RECT  5.670 0.540 5.830 2.460 ;
        RECT  4.890 1.070 5.050 1.350 ;
        RECT  4.890 1.130 5.830 1.290 ;
        RECT  2.930 2.600 5.060 2.760 ;
        RECT  4.900 2.420 5.060 2.760 ;
        RECT  3.890 0.820 4.050 2.760 ;
        RECT  2.930 2.150 3.090 2.760 ;
        RECT  4.900 2.420 5.430 2.580 ;
        RECT  5.270 1.550 5.430 2.580 ;
        RECT  1.890 2.150 3.090 2.310 ;
        RECT  3.710 0.820 4.050 0.980 ;
        RECT  4.530 2.130 4.740 2.440 ;
        RECT  4.530 0.540 4.690 2.440 ;
        RECT  0.100 2.300 1.010 2.460 ;
        RECT  0.850 0.560 1.010 2.460 ;
        RECT  4.210 0.440 4.370 2.060 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  0.850 0.560 2.490 0.720 ;
        RECT  2.330 0.440 4.370 0.600 ;
        RECT  3.270 2.150 3.730 2.310 ;
        RECT  3.570 1.140 3.730 2.310 ;
        RECT  3.350 1.140 3.730 1.300 ;
        RECT  3.350 0.820 3.510 1.300 ;
        RECT  3.230 0.820 3.510 1.040 ;
        RECT  1.290 0.880 1.450 2.120 ;
        RECT  1.290 1.830 3.410 1.990 ;
        RECT  3.250 1.510 3.410 1.990 ;
        RECT  1.290 0.880 1.580 1.100 ;
    END
END DBAHRBEHD

MACRO DBAHRBHHD
    CLASS CORE ;
    FOREIGN DBAHRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.000 2.300 1.650 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 0.900 8.300 2.300 ;
        RECT  7.820 2.100 8.300 2.300 ;
        RECT  7.820 0.900 8.300 1.100 ;
        END
    END QB
    PIN GB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END GB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.370 2.970 1.650 ;
        RECT  2.500 1.000 2.700 1.650 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.850 7.100 2.120 ;
        RECT  6.760 1.840 7.100 2.120 ;
        RECT  6.760 0.850 7.100 1.130 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.980 ;
        RECT  6.180 -0.280 6.460 0.580 ;
        RECT  7.300 -0.280 7.580 0.580 ;
        RECT  8.420 -0.280 8.700 0.580 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.620 2.800 3.480 ;
        RECT  5.240 2.320 5.460 3.480 ;
        RECT  6.180 2.620 6.460 3.480 ;
        RECT  7.260 2.620 7.540 3.480 ;
        RECT  8.380 2.620 8.660 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.760 2.300 7.620 2.460 ;
        RECT  7.460 1.420 7.620 2.460 ;
        RECT  5.760 0.820 5.920 2.460 ;
        RECT  4.890 1.140 5.110 1.420 ;
        RECT  4.890 1.200 5.920 1.360 ;
        RECT  5.700 0.820 5.980 0.980 ;
        RECT  2.970 2.600 5.070 2.760 ;
        RECT  4.910 1.940 5.070 2.760 ;
        RECT  3.930 0.760 4.090 2.760 ;
        RECT  2.970 2.300 3.130 2.760 ;
        RECT  1.930 2.300 3.130 2.460 ;
        RECT  4.910 1.940 5.590 2.100 ;
        RECT  5.370 1.560 5.590 2.100 ;
        RECT  4.560 2.130 4.750 2.440 ;
        RECT  4.570 0.760 4.730 2.440 ;
        RECT  0.100 2.300 1.010 2.460 ;
        RECT  0.850 0.580 1.010 2.460 ;
        RECT  0.100 2.220 0.380 2.460 ;
        RECT  4.250 0.440 4.410 2.070 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.850 0.580 2.490 0.740 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.330 0.440 4.410 0.600 ;
        RECT  3.310 2.240 3.770 2.400 ;
        RECT  3.610 0.940 3.770 2.400 ;
        RECT  3.190 0.940 3.770 1.100 ;
        RECT  3.190 0.820 3.410 1.100 ;
        RECT  1.290 0.900 1.450 2.120 ;
        RECT  1.290 1.920 3.450 2.080 ;
        RECT  3.290 1.480 3.450 2.080 ;
        RECT  1.250 0.900 1.530 1.120 ;
    END
END DBAHRBHHD

MACRO DBFRBEHD
    CLASS CORE ;
    FOREIGN DBFRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 1.280 7.100 1.940 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.840 9.900 2.390 ;
        RECT  9.680 2.110 9.900 2.390 ;
        RECT  9.680 0.840 9.900 1.120 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.280 1.500 1.850 ;
        RECT  1.180 1.440 1.500 1.720 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.640 1.840 8.860 2.120 ;
        RECT  8.640 1.040 9.100 1.240 ;
        RECT  8.900 1.040 9.100 2.040 ;
        RECT  8.640 1.840 9.100 2.040 ;
        RECT  8.640 0.960 8.860 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.240 -0.280 1.520 0.400 ;
        RECT  6.740 -0.280 7.020 0.400 ;
        RECT  7.680 -0.280 7.960 0.400 ;
        RECT  9.100 -0.280 9.380 0.580 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.800 1.660 3.480 ;
        RECT  6.220 2.800 6.500 3.480 ;
        RECT  6.670 2.800 6.950 3.480 ;
        RECT  6.220 2.860 6.950 3.480 ;
        RECT  9.100 2.620 9.380 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.200 2.600 4.280 2.760 ;
        RECT  4.120 2.140 4.280 2.760 ;
        RECT  6.000 2.480 8.450 2.640 ;
        RECT  8.290 0.440 8.450 2.640 ;
        RECT  3.200 0.460 3.360 2.760 ;
        RECT  2.820 2.300 3.360 2.520 ;
        RECT  6.000 2.140 6.160 2.640 ;
        RECT  8.290 2.300 9.480 2.460 ;
        RECT  9.320 1.300 9.480 2.460 ;
        RECT  4.120 2.140 6.160 2.300 ;
        RECT  3.040 0.460 3.360 0.680 ;
        RECT  8.240 0.440 8.520 0.660 ;
        RECT  7.190 2.160 7.950 2.320 ;
        RECT  7.790 0.980 7.950 2.320 ;
        RECT  7.790 1.460 8.110 1.740 ;
        RECT  3.520 2.220 3.850 2.440 ;
        RECT  3.520 0.440 3.680 2.440 ;
        RECT  7.470 0.620 7.630 1.720 ;
        RECT  6.420 0.620 7.630 0.780 ;
        RECT  6.420 0.440 6.580 0.780 ;
        RECT  3.520 0.440 6.580 0.600 ;
        RECT  6.320 1.820 6.480 2.220 ;
        RECT  4.420 1.820 6.480 1.980 ;
        RECT  5.620 1.080 5.780 1.980 ;
        RECT  5.620 1.080 5.940 1.300 ;
        RECT  4.360 1.080 5.940 1.240 ;
        RECT  4.360 0.840 4.520 1.240 ;
        RECT  5.940 1.460 6.260 1.620 ;
        RECT  6.100 0.760 6.260 1.620 ;
        RECT  4.780 0.760 6.260 0.920 ;
        RECT  5.620 2.460 5.840 2.740 ;
        RECT  4.700 2.460 5.840 2.620 ;
        RECT  3.840 1.400 4.220 1.980 ;
        RECT  3.840 1.400 5.310 1.560 ;
        RECT  3.840 0.840 4.000 1.980 ;
        RECT  0.600 1.710 0.760 2.180 ;
        RECT  2.880 0.880 3.040 2.080 ;
        RECT  0.580 0.440 0.740 1.870 ;
        RECT  2.720 0.520 2.880 1.040 ;
        RECT  0.580 0.560 1.840 0.720 ;
        RECT  1.680 0.520 2.880 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.000 2.530 2.660 2.690 ;
        RECT  2.000 0.840 2.160 2.690 ;
        RECT  2.000 0.840 2.550 1.120 ;
        RECT  0.900 2.380 1.840 2.540 ;
        RECT  1.680 0.920 1.840 2.540 ;
        RECT  0.900 0.920 1.840 1.080 ;
    END
END DBFRBEHD

MACRO DBFRBHHD
    CLASS CORE ;
    FOREIGN DBFRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.790 10.700 2.360 ;
        RECT  10.360 2.080 10.700 2.360 ;
        RECT  10.360 0.820 10.700 1.100 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.200 1.500 1.740 ;
        RECT  1.260 1.440 1.500 1.720 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.610 9.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.580 -0.280 1.860 0.400 ;
        RECT  6.760 -0.280 7.040 0.400 ;
        RECT  8.740 -0.280 9.020 0.580 ;
        RECT  9.780 -0.280 10.060 0.580 ;
        RECT  10.820 -0.280 11.100 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.580 2.800 1.860 3.480 ;
        RECT  6.820 2.740 7.160 3.480 ;
        RECT  7.840 2.620 8.120 3.480 ;
        RECT  8.740 2.620 9.020 3.480 ;
        RECT  9.780 2.620 10.060 3.480 ;
        RECT  10.820 2.620 11.100 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.170 2.600 6.660 2.760 ;
        RECT  6.500 2.420 6.660 2.760 ;
        RECT  3.170 0.460 3.330 2.760 ;
        RECT  6.500 2.420 7.630 2.580 ;
        RECT  2.790 2.300 3.330 2.520 ;
        RECT  10.040 1.420 10.200 2.460 ;
        RECT  7.470 2.300 10.200 2.460 ;
        RECT  8.240 1.940 8.520 2.460 ;
        RECT  8.360 0.950 8.520 2.460 ;
        RECT  8.240 0.950 8.520 1.230 ;
        RECT  3.010 0.460 3.330 0.680 ;
        RECT  7.280 1.980 8.020 2.140 ;
        RECT  7.860 0.630 8.020 2.140 ;
        RECT  7.860 1.460 8.200 1.740 ;
        RECT  7.700 0.630 8.020 0.910 ;
        RECT  3.490 2.220 3.820 2.440 ;
        RECT  3.490 0.440 3.650 2.440 ;
        RECT  7.360 1.400 7.680 1.680 ;
        RECT  7.360 0.560 7.520 1.680 ;
        RECT  6.370 0.560 7.520 0.720 ;
        RECT  3.490 0.440 6.530 0.600 ;
        RECT  4.760 2.280 6.340 2.440 ;
        RECT  6.180 1.460 6.340 2.440 ;
        RECT  5.790 1.460 6.340 1.620 ;
        RECT  6.050 0.760 6.210 1.620 ;
        RECT  4.710 0.760 6.210 0.920 ;
        RECT  5.070 1.960 6.020 2.120 ;
        RECT  5.740 1.900 6.020 2.120 ;
        RECT  4.390 1.820 5.230 1.980 ;
        RECT  5.070 1.080 5.230 2.120 ;
        RECT  5.610 1.080 5.890 1.300 ;
        RECT  4.330 1.080 5.890 1.240 ;
        RECT  4.330 0.840 4.490 1.240 ;
        RECT  3.810 1.400 4.190 1.980 ;
        RECT  3.810 1.400 4.900 1.560 ;
        RECT  3.810 0.840 3.970 1.980 ;
        RECT  0.600 2.480 2.630 2.640 ;
        RECT  2.470 1.980 2.630 2.640 ;
        RECT  0.600 1.680 0.760 2.640 ;
        RECT  2.470 1.980 3.010 2.140 ;
        RECT  2.850 0.840 3.010 2.140 ;
        RECT  0.580 0.440 0.740 1.840 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.140 1.640 2.300 2.290 ;
        RECT  2.200 1.580 2.640 1.800 ;
        RECT  2.200 0.550 2.360 1.800 ;
        RECT  2.200 0.550 2.720 0.710 ;
        RECT  0.980 2.160 1.950 2.320 ;
        RECT  1.790 0.880 1.950 2.320 ;
        RECT  0.980 0.880 1.950 1.040 ;
    END
END DBFRBHHD

MACRO DBFRSBEHD
    CLASS CORE ;
    FOREIGN DBFRSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.170 0.840 7.500 1.340 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.480 1.840 10.700 2.120 ;
        RECT  10.500 0.920 10.700 2.160 ;
        RECT  10.480 0.960 10.700 1.240 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.190 1.420 1.500 1.700 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.090 0.700 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.960 9.900 2.120 ;
        RECT  9.380 1.840 9.900 2.120 ;
        RECT  9.380 0.960 9.900 1.240 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.420 8.310 1.700 ;
        RECT  8.100 1.420 8.300 1.960 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.270 -0.280 1.550 0.400 ;
        RECT  5.550 -0.280 5.830 0.620 ;
        RECT  6.950 -0.280 7.230 0.620 ;
        RECT  8.170 -0.280 8.450 0.620 ;
        RECT  9.900 -0.280 10.180 0.580 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 2.800 1.680 3.480 ;
        RECT  5.050 2.800 5.330 3.480 ;
        RECT  6.710 2.480 6.970 3.480 ;
        RECT  7.770 2.800 8.050 3.480 ;
        RECT  8.790 2.800 9.070 3.480 ;
        RECT  9.900 2.620 10.180 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.670 2.800 0.950 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.010 2.600 4.240 2.760 ;
        RECT  4.080 2.160 4.240 2.760 ;
        RECT  3.010 0.460 3.170 2.760 ;
        RECT  2.690 2.300 3.170 2.520 ;
        RECT  9.000 2.280 10.280 2.440 ;
        RECT  10.120 1.300 10.280 2.440 ;
        RECT  4.080 2.160 9.160 2.320 ;
        RECT  9.000 0.440 9.160 2.440 ;
        RECT  9.000 0.440 9.290 0.750 ;
        RECT  2.850 0.460 3.170 0.680 ;
        RECT  8.630 1.090 8.790 1.460 ;
        RECT  8.520 1.090 8.790 1.250 ;
        RECT  7.830 0.940 8.680 1.100 ;
        RECT  8.300 2.480 8.630 2.740 ;
        RECT  7.130 2.480 8.630 2.640 ;
        RECT  3.640 2.280 3.920 2.440 ;
        RECT  3.680 1.840 3.840 2.440 ;
        RECT  3.680 1.840 4.570 2.000 ;
        RECT  4.410 1.060 4.570 2.000 ;
        RECT  7.570 1.500 7.730 1.920 ;
        RECT  4.410 1.500 7.730 1.660 ;
        RECT  3.990 1.060 4.570 1.220 ;
        RECT  3.990 0.600 4.150 1.220 ;
        RECT  3.370 0.600 4.150 0.760 ;
        RECT  3.370 0.460 3.710 0.760 ;
        RECT  4.730 1.820 7.410 1.980 ;
        RECT  4.400 2.480 6.550 2.640 ;
        RECT  4.840 1.180 6.290 1.340 ;
        RECT  6.130 0.700 6.290 1.340 ;
        RECT  4.840 0.880 5.000 1.340 ;
        RECT  4.730 0.880 5.000 1.160 ;
        RECT  5.160 0.780 5.970 1.020 ;
        RECT  5.160 0.460 5.320 1.020 ;
        RECT  4.340 0.460 5.320 0.620 ;
        RECT  3.330 0.940 3.490 2.080 ;
        RECT  3.330 1.380 4.250 1.660 ;
        RECT  3.330 0.940 3.690 1.100 ;
        RECT  0.160 0.450 0.320 2.700 ;
        RECT  0.160 2.480 2.500 2.640 ;
        RECT  2.340 1.960 2.500 2.640 ;
        RECT  2.340 1.960 2.850 2.120 ;
        RECT  2.690 0.840 2.850 2.120 ;
        RECT  0.100 0.450 0.380 0.710 ;
        RECT  2.020 0.520 2.180 2.310 ;
        RECT  2.020 1.540 2.380 1.800 ;
        RECT  2.020 0.520 2.670 0.680 ;
        RECT  0.920 2.120 1.820 2.280 ;
        RECT  1.660 0.920 1.820 2.280 ;
        RECT  1.660 1.410 1.860 1.800 ;
        RECT  0.920 0.920 1.820 1.080 ;
    END
END DBFRSBEHD

MACRO DBFRSBHHD
    CLASS CORE ;
    FOREIGN DBFRSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 1.360 7.500 1.990 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.920 11.500 2.160 ;
        RECT  11.160 1.840 11.500 2.160 ;
        RECT  11.160 0.920 11.500 1.240 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.190 1.420 1.500 1.700 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.090 0.700 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.060 0.960 10.340 1.240 ;
        RECT  10.060 1.840 10.340 2.120 ;
        RECT  10.100 0.960 10.300 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.270 8.700 1.960 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 -0.280 1.680 0.400 ;
        RECT  5.530 -0.280 5.750 0.680 ;
        RECT  7.050 -0.280 7.330 0.620 ;
        RECT  8.270 -0.280 8.550 0.620 ;
        RECT  9.500 -0.280 9.780 0.400 ;
        RECT  10.580 -0.280 10.860 0.580 ;
        RECT  11.620 -0.280 11.900 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 2.800 1.680 3.480 ;
        RECT  4.980 2.800 5.260 3.480 ;
        RECT  6.340 2.800 6.620 3.480 ;
        RECT  7.080 2.800 7.360 3.480 ;
        RECT  8.460 2.800 8.740 3.480 ;
        RECT  9.540 2.600 9.820 3.480 ;
        RECT  10.580 2.620 10.860 3.480 ;
        RECT  11.620 2.620 11.900 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.020 2.480 9.380 2.760 ;
        RECT  9.220 2.280 9.380 2.760 ;
        RECT  2.680 2.600 4.170 2.760 ;
        RECT  4.010 2.160 4.170 2.760 ;
        RECT  6.440 2.480 9.380 2.640 ;
        RECT  2.680 2.300 3.100 2.760 ;
        RECT  2.940 0.460 3.100 2.760 ;
        RECT  6.440 2.160 6.600 2.640 ;
        RECT  9.220 2.280 11.000 2.440 ;
        RECT  10.840 1.300 11.000 2.440 ;
        RECT  4.010 2.160 6.600 2.320 ;
        RECT  9.410 0.780 9.570 2.440 ;
        RECT  9.170 0.780 9.570 0.940 ;
        RECT  9.170 0.660 9.390 0.940 ;
        RECT  2.780 0.460 3.100 0.680 ;
        RECT  7.640 2.160 9.060 2.320 ;
        RECT  8.900 1.470 9.060 2.320 ;
        RECT  8.160 1.220 8.320 2.320 ;
        RECT  8.900 1.470 9.240 1.750 ;
        RECT  7.990 1.220 8.320 1.500 ;
        RECT  3.570 2.280 3.850 2.440 ;
        RECT  3.610 1.840 3.770 2.440 ;
        RECT  3.610 1.840 4.500 2.000 ;
        RECT  4.340 1.060 4.500 2.000 ;
        RECT  7.660 1.660 8.000 1.940 ;
        RECT  4.340 1.500 6.820 1.660 ;
        RECT  6.660 0.880 6.820 1.660 ;
        RECT  7.660 0.880 7.820 1.940 ;
        RECT  3.920 1.060 4.500 1.220 ;
        RECT  3.920 0.600 4.080 1.220 ;
        RECT  6.660 0.880 7.820 1.040 ;
        RECT  3.300 0.600 4.080 0.760 ;
        RECT  3.300 0.460 3.640 0.760 ;
        RECT  6.760 2.160 7.100 2.320 ;
        RECT  6.760 1.820 6.920 2.320 ;
        RECT  4.660 1.820 6.920 1.980 ;
        RECT  5.090 0.840 6.070 1.000 ;
        RECT  5.910 0.560 6.070 1.000 ;
        RECT  5.090 0.460 5.250 1.000 ;
        RECT  5.910 0.560 6.630 0.720 ;
        RECT  4.270 0.460 5.250 0.620 ;
        RECT  4.770 1.180 6.450 1.340 ;
        RECT  6.230 0.880 6.450 1.340 ;
        RECT  4.770 0.880 4.930 1.340 ;
        RECT  4.660 0.880 4.930 1.160 ;
        RECT  4.330 2.480 6.280 2.640 ;
        RECT  3.260 0.940 3.420 2.080 ;
        RECT  3.260 1.380 4.180 1.660 ;
        RECT  3.260 0.940 3.620 1.100 ;
        RECT  0.100 2.380 0.380 2.660 ;
        RECT  0.100 2.480 2.500 2.640 ;
        RECT  2.340 1.980 2.500 2.640 ;
        RECT  0.160 0.480 0.320 2.660 ;
        RECT  2.340 1.980 2.780 2.140 ;
        RECT  2.620 0.840 2.780 2.140 ;
        RECT  0.100 0.480 0.380 0.700 ;
        RECT  2.020 0.530 2.180 2.280 ;
        RECT  2.020 1.580 2.420 1.800 ;
        RECT  2.020 0.530 2.520 0.690 ;
        RECT  0.920 2.160 1.840 2.320 ;
        RECT  1.680 0.880 1.840 2.320 ;
        RECT  0.920 0.880 1.840 1.040 ;
    END
END DBFRSBHHD

MACRO DBZRBEHD
    CLASS CORE ;
    FOREIGN DBZRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.280 9.100 1.940 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 0.840 11.900 2.390 ;
        RECT  11.680 2.110 11.900 2.390 ;
        RECT  11.680 0.840 11.900 1.120 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.200 3.500 1.740 ;
        RECT  3.260 1.440 3.500 1.720 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.000 11.100 2.080 ;
        RECT  10.580 1.880 11.100 2.080 ;
        RECT  10.580 1.000 11.100 1.200 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.570 -0.280 3.850 0.400 ;
        RECT  8.710 -0.280 8.990 0.400 ;
        RECT  9.680 -0.280 9.960 0.400 ;
        RECT  11.100 -0.280 11.380 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.530 2.800 3.810 3.480 ;
        RECT  8.190 2.800 8.920 3.480 ;
        RECT  9.760 2.800 10.040 3.480 ;
        RECT  11.100 2.620 11.380 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.170 2.600 6.250 2.760 ;
        RECT  6.090 2.140 6.250 2.760 ;
        RECT  7.970 2.480 10.460 2.640 ;
        RECT  10.260 2.300 10.460 2.640 ;
        RECT  5.170 0.460 5.330 2.760 ;
        RECT  4.790 2.300 5.330 2.520 ;
        RECT  7.970 2.140 8.130 2.640 ;
        RECT  10.260 2.300 11.480 2.460 ;
        RECT  11.320 1.300 11.480 2.460 ;
        RECT  6.090 2.140 8.130 2.300 ;
        RECT  10.260 0.440 10.420 2.640 ;
        RECT  10.260 0.440 10.460 0.720 ;
        RECT  5.010 0.460 5.330 0.680 ;
        RECT  9.160 2.160 9.920 2.320 ;
        RECT  9.760 0.980 9.920 2.320 ;
        RECT  9.760 1.460 10.080 1.740 ;
        RECT  5.490 2.220 5.820 2.440 ;
        RECT  5.490 0.440 5.650 2.440 ;
        RECT  9.440 0.620 9.600 1.720 ;
        RECT  8.390 0.620 9.600 0.780 ;
        RECT  8.390 0.440 8.550 0.780 ;
        RECT  5.490 0.440 8.550 0.600 ;
        RECT  8.290 1.820 8.450 2.220 ;
        RECT  6.390 1.820 8.450 1.980 ;
        RECT  7.590 1.080 7.750 1.980 ;
        RECT  7.590 1.080 7.910 1.300 ;
        RECT  6.330 1.080 7.910 1.240 ;
        RECT  6.330 0.840 6.490 1.240 ;
        RECT  7.910 1.460 8.230 1.620 ;
        RECT  8.070 0.760 8.230 1.620 ;
        RECT  6.750 0.760 8.230 0.920 ;
        RECT  7.590 2.460 7.810 2.740 ;
        RECT  6.670 2.460 7.810 2.620 ;
        RECT  5.810 1.400 6.190 1.980 ;
        RECT  5.810 1.400 7.280 1.560 ;
        RECT  5.810 0.840 5.970 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.470 1.980 4.630 2.640 ;
        RECT  2.200 2.480 4.630 2.640 ;
        RECT  4.470 1.980 5.010 2.140 ;
        RECT  4.850 0.840 5.010 2.140 ;
        RECT  1.620 0.560 2.360 0.720 ;
        RECT  4.150 1.640 4.310 2.310 ;
        RECT  4.190 1.580 4.590 1.800 ;
        RECT  4.190 0.560 4.350 1.800 ;
        RECT  4.190 0.560 4.690 0.720 ;
        RECT  2.930 2.160 3.900 2.320 ;
        RECT  3.740 0.880 3.900 2.320 ;
        RECT  2.930 0.880 3.900 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.790 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END DBZRBEHD

MACRO DBZRBHHD
    CLASS CORE ;
    FOREIGN DBZRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.400 8.760 1.680 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 0.790 12.700 2.360 ;
        RECT  12.360 2.080 12.700 2.360 ;
        RECT  12.360 0.820 12.700 1.100 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.200 3.500 1.740 ;
        RECT  3.260 1.260 3.500 1.540 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.610 11.500 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.420 -0.280 3.700 0.400 ;
        RECT  8.690 -0.280 8.970 0.400 ;
        RECT  10.740 -0.280 11.020 0.580 ;
        RECT  11.780 -0.280 12.060 0.580 ;
        RECT  12.820 -0.280 13.100 0.580 ;
        RECT  0.000 -0.280 13.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.420 2.800 3.700 3.480 ;
        RECT  8.750 2.740 9.090 3.480 ;
        RECT  9.770 2.620 10.050 3.480 ;
        RECT  10.740 2.620 11.020 3.480 ;
        RECT  11.780 2.620 12.060 3.480 ;
        RECT  12.820 2.620 13.100 3.480 ;
        RECT  0.000 2.920 13.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.100 2.600 8.590 2.760 ;
        RECT  8.430 2.420 8.590 2.760 ;
        RECT  5.100 0.460 5.260 2.760 ;
        RECT  8.430 2.420 9.560 2.580 ;
        RECT  4.720 2.300 5.260 2.520 ;
        RECT  12.040 1.420 12.200 2.460 ;
        RECT  9.400 2.300 12.200 2.460 ;
        RECT  10.240 1.940 10.460 2.460 ;
        RECT  10.300 0.960 10.460 2.460 ;
        RECT  10.240 0.960 10.460 1.240 ;
        RECT  4.940 0.460 5.260 0.680 ;
        RECT  9.310 1.860 9.930 2.140 ;
        RECT  9.770 0.480 9.930 2.140 ;
        RECT  9.770 1.460 10.130 1.740 ;
        RECT  9.630 0.480 9.930 0.760 ;
        RECT  5.420 2.220 5.750 2.440 ;
        RECT  5.420 0.440 5.580 2.440 ;
        RECT  9.290 1.400 9.610 1.680 ;
        RECT  9.290 0.560 9.450 1.680 ;
        RECT  8.300 0.560 9.450 0.720 ;
        RECT  5.420 0.440 8.460 0.600 ;
        RECT  6.690 2.280 8.270 2.440 ;
        RECT  8.110 1.460 8.270 2.440 ;
        RECT  7.720 1.460 8.270 1.620 ;
        RECT  7.980 0.760 8.140 1.620 ;
        RECT  6.640 0.760 8.140 0.920 ;
        RECT  7.000 1.960 7.950 2.120 ;
        RECT  7.670 1.900 7.950 2.120 ;
        RECT  6.320 1.820 7.160 1.980 ;
        RECT  7.000 1.080 7.160 2.120 ;
        RECT  7.540 1.080 7.820 1.300 ;
        RECT  6.260 1.080 7.820 1.240 ;
        RECT  6.260 0.840 6.420 1.240 ;
        RECT  5.740 1.400 6.120 1.980 ;
        RECT  5.740 1.400 6.830 1.560 ;
        RECT  5.740 0.840 5.900 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.400 1.980 4.560 2.640 ;
        RECT  2.200 2.480 4.560 2.640 ;
        RECT  4.400 1.980 4.940 2.140 ;
        RECT  4.780 0.840 4.940 2.140 ;
        RECT  1.610 0.560 2.360 0.720 ;
        RECT  4.080 0.520 4.240 2.300 ;
        RECT  4.080 1.580 4.520 1.800 ;
        RECT  4.080 0.520 4.750 0.680 ;
        RECT  2.820 2.160 3.900 2.320 ;
        RECT  3.740 0.880 3.900 2.320 ;
        RECT  2.820 0.880 3.900 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END DBZRBHHD

MACRO DBZRSBEHD
    CLASS CORE ;
    FOREIGN DBZRSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.800 0.840 9.100 1.340 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.420 2.300 1.990 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.080 1.840 12.300 2.120 ;
        RECT  12.100 0.920 12.300 2.160 ;
        RECT  12.080 0.960 12.300 1.240 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.100 1.960 ;
        RECT  2.890 1.420 3.100 1.700 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.960 11.260 1.240 ;
        RECT  10.900 1.840 11.260 2.120 ;
        RECT  10.900 0.960 11.100 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 1.420 9.940 1.700 ;
        RECT  9.700 1.420 9.900 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.400 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.500 -0.280 3.220 0.400 ;
        RECT  7.180 -0.280 7.460 0.620 ;
        RECT  8.580 -0.280 8.860 0.620 ;
        RECT  9.800 -0.280 10.080 0.620 ;
        RECT  11.500 -0.280 11.780 0.580 ;
        RECT  0.000 -0.280 12.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 2.800 2.620 3.480 ;
        RECT  3.100 2.800 3.380 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  8.240 2.800 8.520 3.480 ;
        RECT  9.400 2.800 9.680 3.480 ;
        RECT  10.420 2.800 10.700 3.480 ;
        RECT  11.500 2.620 11.780 3.480 ;
        RECT  0.000 2.920 12.400 3.480 ;
        RECT  0.520 2.620 0.800 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.380 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  4.380 2.300 4.800 2.760 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  10.580 2.280 11.880 2.440 ;
        RECT  11.720 1.300 11.880 2.440 ;
        RECT  5.710 2.160 10.740 2.320 ;
        RECT  10.580 0.440 10.740 2.440 ;
        RECT  10.580 0.440 10.920 0.750 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  10.260 0.940 10.420 1.460 ;
        RECT  9.460 0.940 10.420 1.100 ;
        RECT  9.930 2.480 10.260 2.740 ;
        RECT  8.760 2.480 10.260 2.640 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  9.200 1.500 9.360 1.920 ;
        RECT  6.040 1.500 9.360 1.660 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  6.360 1.820 9.040 1.980 ;
        RECT  6.030 2.480 8.180 2.640 ;
        RECT  6.470 1.180 7.920 1.340 ;
        RECT  7.760 0.700 7.920 1.340 ;
        RECT  6.470 0.880 6.630 1.340 ;
        RECT  6.360 0.880 6.630 1.160 ;
        RECT  6.790 0.780 7.600 1.000 ;
        RECT  6.790 0.460 6.950 1.000 ;
        RECT  5.970 0.460 6.950 0.620 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  2.280 2.480 4.220 2.640 ;
        RECT  4.060 1.960 4.220 2.640 ;
        RECT  2.280 2.220 2.440 2.640 ;
        RECT  1.320 2.220 2.440 2.380 ;
        RECT  1.720 0.460 1.880 2.380 ;
        RECT  4.060 1.960 4.480 2.120 ;
        RECT  4.320 0.840 4.480 2.120 ;
        RECT  1.620 0.460 1.900 0.680 ;
        RECT  3.720 0.520 3.880 2.320 ;
        RECT  3.720 1.640 4.120 1.800 ;
        RECT  3.720 0.520 4.230 0.680 ;
        RECT  2.620 2.160 3.540 2.320 ;
        RECT  3.380 0.940 3.540 2.320 ;
        RECT  2.620 0.940 3.540 1.100 ;
        RECT  0.980 2.600 1.920 2.760 ;
        RECT  0.980 2.200 1.140 2.760 ;
        RECT  0.880 1.060 1.040 2.360 ;
        RECT  0.080 1.060 0.240 2.320 ;
        RECT  0.080 2.000 0.320 2.280 ;
        RECT  0.080 1.060 1.040 1.220 ;
        RECT  0.100 0.740 0.380 1.220 ;
    END
END DBZRSBEHD

MACRO DBZRSBHHD
    CLASS CORE ;
    FOREIGN DBZRSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 1.510 9.500 2.140 ;
        END
    END RB
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.420 2.700 1.990 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 0.920 13.500 2.160 ;
        RECT  13.160 1.840 13.500 2.160 ;
        RECT  13.160 0.920 13.500 1.240 ;
        END
    END QB
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.420 3.500 1.960 ;
        RECT  3.180 1.420 3.500 1.700 ;
        END
    END CKB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.060 0.960 12.340 1.240 ;
        RECT  12.060 1.840 12.340 2.120 ;
        RECT  12.100 0.960 12.300 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.350 10.700 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.280 2.800 0.400 ;
        RECT  3.220 -0.280 3.500 0.400 ;
        RECT  7.510 -0.280 7.730 0.680 ;
        RECT  9.030 -0.280 9.310 0.620 ;
        RECT  10.320 -0.280 10.600 0.620 ;
        RECT  11.500 -0.280 11.780 0.400 ;
        RECT  12.580 -0.280 12.860 0.580 ;
        RECT  13.620 -0.280 13.900 0.580 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.380 2.800 3.660 3.480 ;
        RECT  6.960 2.800 7.240 3.480 ;
        RECT  8.380 2.800 8.660 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  10.380 2.800 10.660 3.480 ;
        RECT  11.500 2.800 11.780 3.480 ;
        RECT  12.580 2.620 12.860 3.480 ;
        RECT  13.620 2.620 13.900 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 6.150 2.760 ;
        RECT  5.990 2.160 6.150 2.760 ;
        RECT  8.480 2.480 12.350 2.640 ;
        RECT  12.190 2.280 12.350 2.640 ;
        RECT  4.640 2.300 5.080 2.760 ;
        RECT  4.920 0.460 5.080 2.760 ;
        RECT  11.720 0.900 11.880 2.640 ;
        RECT  8.480 2.160 8.640 2.640 ;
        RECT  12.190 2.280 13.000 2.440 ;
        RECT  12.840 1.300 13.000 2.440 ;
        RECT  5.990 2.160 8.640 2.320 ;
        RECT  11.220 0.900 11.880 1.060 ;
        RECT  11.220 0.750 11.440 1.060 ;
        RECT  4.760 0.460 5.080 0.680 ;
        RECT  9.740 2.160 11.480 2.320 ;
        RECT  11.320 1.240 11.480 2.320 ;
        RECT  10.880 1.240 11.480 1.400 ;
        RECT  10.880 0.780 11.040 1.400 ;
        RECT  9.980 0.780 10.230 1.150 ;
        RECT  9.980 0.780 11.040 0.940 ;
        RECT  5.550 2.280 5.830 2.440 ;
        RECT  5.590 1.840 5.750 2.440 ;
        RECT  5.590 1.840 6.480 2.000 ;
        RECT  6.320 1.060 6.480 2.000 ;
        RECT  10.060 1.310 10.220 1.940 ;
        RECT  6.320 1.500 8.800 1.660 ;
        RECT  8.640 0.880 8.800 1.660 ;
        RECT  9.660 1.310 10.220 1.470 ;
        RECT  9.660 0.880 9.820 1.470 ;
        RECT  5.900 1.060 6.480 1.220 ;
        RECT  5.900 0.600 6.060 1.220 ;
        RECT  8.640 0.880 9.820 1.040 ;
        RECT  5.280 0.600 6.060 0.760 ;
        RECT  5.280 0.460 5.620 0.760 ;
        RECT  8.800 2.100 9.140 2.320 ;
        RECT  8.800 1.820 8.960 2.320 ;
        RECT  6.640 1.820 8.960 1.980 ;
        RECT  7.070 0.840 8.050 1.000 ;
        RECT  7.890 0.560 8.050 1.000 ;
        RECT  7.070 0.460 7.230 1.000 ;
        RECT  7.890 0.560 8.610 0.720 ;
        RECT  6.250 0.460 7.230 0.620 ;
        RECT  6.750 1.180 8.430 1.340 ;
        RECT  8.210 0.880 8.430 1.340 ;
        RECT  6.750 0.880 6.910 1.340 ;
        RECT  6.640 0.880 6.910 1.160 ;
        RECT  6.310 2.480 8.320 2.640 ;
        RECT  5.240 0.940 5.400 2.080 ;
        RECT  5.240 1.380 6.160 1.660 ;
        RECT  5.240 0.940 5.600 1.100 ;
        RECT  1.480 2.520 2.340 2.680 ;
        RECT  2.180 0.740 2.340 2.680 ;
        RECT  4.320 1.960 4.480 2.640 ;
        RECT  2.180 2.480 4.480 2.640 ;
        RECT  4.320 1.960 4.760 2.120 ;
        RECT  4.600 0.840 4.760 2.120 ;
        RECT  1.600 0.740 2.340 0.900 ;
        RECT  4.000 0.520 4.160 2.320 ;
        RECT  4.000 1.640 4.400 1.800 ;
        RECT  4.000 0.520 4.500 0.680 ;
        RECT  2.900 2.160 3.820 2.320 ;
        RECT  3.660 0.880 3.820 2.320 ;
        RECT  2.900 0.880 3.820 1.040 ;
        RECT  0.900 2.200 2.020 2.360 ;
        RECT  1.860 1.420 2.020 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END DBZRSBHHD

MACRO DELAKHD
    CLASS CORE ;
    FOREIGN DELAKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.760 6.780 1.080 ;
        RECT  7.550 0.760 7.830 1.080 ;
        RECT  7.700 0.920 7.900 2.280 ;
        RECT  8.600 0.760 8.880 1.080 ;
        RECT  6.500 0.920 8.880 1.080 ;
        RECT  6.560 2.120 8.920 2.280 ;
        RECT  6.560 2.060 6.720 2.340 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.280 1.230 1.560 ;
        RECT  0.900 0.920 1.100 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.720 -0.280 3.000 0.860 ;
        RECT  5.500 -0.280 5.780 0.860 ;
        RECT  7.020 -0.280 7.300 0.760 ;
        RECT  8.070 -0.280 8.350 0.760 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.160 -0.280 0.320 1.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.520 0.980 0.680 2.320 ;
        RECT  0.100 2.160 0.680 2.320 ;
        RECT  2.720 2.400 3.000 3.480 ;
        RECT  5.500 2.400 5.780 3.480 ;
        RECT  7.020 2.620 7.300 3.480 ;
        RECT  8.070 2.620 8.350 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.120 2.160 0.280 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.080 0.640 6.240 2.480 ;
        RECT  6.080 1.520 6.960 1.680 ;
        RECT  4.300 2.040 5.680 2.200 ;
        RECT  5.520 1.120 5.680 2.200 ;
        RECT  5.520 1.430 5.900 1.710 ;
        RECT  4.360 1.120 5.680 1.280 ;
        RECT  4.360 0.640 4.520 1.280 ;
        RECT  3.880 0.640 4.040 2.480 ;
        RECT  3.880 1.520 4.920 1.680 ;
        RECT  1.720 2.040 2.900 2.200 ;
        RECT  2.740 1.120 2.900 2.200 ;
        RECT  2.740 1.430 3.280 1.710 ;
        RECT  1.780 1.120 2.900 1.280 ;
        RECT  1.780 0.640 1.940 1.280 ;
        RECT  1.290 2.240 1.560 2.520 ;
        RECT  1.400 0.640 1.560 2.520 ;
        RECT  1.400 1.520 2.340 1.680 ;
        RECT  1.300 0.640 1.560 0.920 ;
    END
END DELAKHD

MACRO DELBKHD
    CLASS CORE ;
    FOREIGN DELBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.760 6.780 1.080 ;
        RECT  7.550 0.760 7.830 1.080 ;
        RECT  7.700 0.920 7.900 2.280 ;
        RECT  8.600 0.760 8.880 1.080 ;
        RECT  6.500 0.920 8.880 1.080 ;
        RECT  6.560 2.120 8.920 2.280 ;
        RECT  6.560 2.060 6.720 2.340 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.280 1.230 1.560 ;
        RECT  0.900 0.920 1.100 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.720 -0.280 3.000 0.860 ;
        RECT  5.500 -0.280 5.780 0.860 ;
        RECT  7.020 -0.280 7.300 0.760 ;
        RECT  8.070 -0.280 8.350 0.760 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.160 -0.280 0.320 1.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.520 0.980 0.680 2.320 ;
        RECT  0.100 2.160 0.680 2.320 ;
        RECT  2.720 2.400 3.000 3.480 ;
        RECT  5.500 2.400 5.780 3.480 ;
        RECT  7.020 2.620 7.300 3.480 ;
        RECT  8.070 2.620 8.350 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.120 2.160 0.280 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.080 0.640 6.240 2.480 ;
        RECT  6.080 1.520 6.960 1.680 ;
        RECT  4.300 2.040 5.680 2.200 ;
        RECT  5.520 1.120 5.680 2.200 ;
        RECT  5.520 1.430 5.900 1.710 ;
        RECT  4.360 1.120 5.680 1.280 ;
        RECT  4.360 0.640 4.520 1.280 ;
        RECT  3.880 0.640 4.040 2.480 ;
        RECT  3.880 1.520 4.920 1.680 ;
        RECT  1.720 2.040 2.900 2.200 ;
        RECT  2.740 1.120 2.900 2.200 ;
        RECT  2.740 1.430 3.280 1.710 ;
        RECT  1.780 1.120 2.900 1.280 ;
        RECT  1.780 0.640 1.940 1.280 ;
        RECT  1.290 2.240 1.560 2.520 ;
        RECT  1.400 0.640 1.560 2.520 ;
        RECT  1.400 1.520 2.340 1.680 ;
        RECT  1.300 0.640 1.560 0.920 ;
    END
END DELBKHD

MACRO DELCKHD
    CLASS CORE ;
    FOREIGN DELCKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.760 6.780 1.080 ;
        RECT  7.550 0.760 7.830 1.080 ;
        RECT  7.700 0.920 7.900 2.280 ;
        RECT  8.600 0.760 8.880 1.080 ;
        RECT  6.500 0.920 8.880 1.080 ;
        RECT  6.560 2.120 8.920 2.280 ;
        RECT  6.560 2.060 6.720 2.340 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.280 1.230 1.560 ;
        RECT  0.900 0.920 1.100 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.720 -0.280 3.000 0.860 ;
        RECT  5.500 -0.280 5.780 0.860 ;
        RECT  7.020 -0.280 7.300 0.760 ;
        RECT  8.070 -0.280 8.350 0.760 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.160 -0.280 0.320 1.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.520 0.980 0.680 2.320 ;
        RECT  0.100 2.160 0.680 2.320 ;
        RECT  2.720 2.400 3.000 3.480 ;
        RECT  5.500 2.400 5.780 3.480 ;
        RECT  7.020 2.620 7.300 3.480 ;
        RECT  8.070 2.620 8.350 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.120 2.160 0.280 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.080 0.640 6.240 2.480 ;
        RECT  6.080 1.520 6.960 1.680 ;
        RECT  4.300 2.040 5.680 2.200 ;
        RECT  5.520 1.120 5.680 2.200 ;
        RECT  5.520 1.430 5.900 1.710 ;
        RECT  4.360 1.120 5.680 1.280 ;
        RECT  4.360 0.640 4.520 1.280 ;
        RECT  3.880 0.640 4.040 2.480 ;
        RECT  3.880 1.520 4.920 1.680 ;
        RECT  1.720 2.040 2.900 2.200 ;
        RECT  2.740 1.120 2.900 2.200 ;
        RECT  2.740 1.430 3.280 1.710 ;
        RECT  1.780 1.120 2.900 1.280 ;
        RECT  1.780 0.640 1.940 1.280 ;
        RECT  1.290 2.240 1.560 2.520 ;
        RECT  1.400 0.640 1.560 2.520 ;
        RECT  1.400 1.520 2.340 1.680 ;
        RECT  1.300 0.640 1.560 0.920 ;
    END
END DELCKHD

MACRO DELDKHD
    CLASS CORE ;
    FOREIGN DELDKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.760 6.780 1.080 ;
        RECT  7.550 0.760 7.830 1.080 ;
        RECT  7.700 0.920 7.900 2.280 ;
        RECT  8.600 0.760 8.880 1.080 ;
        RECT  6.500 0.920 8.880 1.080 ;
        RECT  6.560 2.120 8.920 2.280 ;
        RECT  6.560 2.060 6.720 2.340 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.280 1.230 1.560 ;
        RECT  0.900 0.920 1.100 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.720 -0.280 3.000 0.860 ;
        RECT  5.500 -0.280 5.780 0.860 ;
        RECT  7.020 -0.280 7.300 0.760 ;
        RECT  8.070 -0.280 8.350 0.760 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.160 -0.280 0.320 1.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.520 0.980 0.680 2.320 ;
        RECT  0.100 2.160 0.680 2.320 ;
        RECT  2.720 2.400 3.000 3.480 ;
        RECT  5.500 2.400 5.780 3.480 ;
        RECT  7.020 2.620 7.300 3.480 ;
        RECT  8.070 2.620 8.350 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.120 2.160 0.280 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.080 0.640 6.240 2.480 ;
        RECT  6.080 1.520 6.960 1.680 ;
        RECT  4.300 2.040 5.680 2.200 ;
        RECT  5.520 1.120 5.680 2.200 ;
        RECT  5.520 1.430 5.900 1.710 ;
        RECT  4.360 1.120 5.680 1.280 ;
        RECT  4.360 0.640 4.520 1.280 ;
        RECT  3.880 0.640 4.040 2.480 ;
        RECT  3.880 1.520 4.920 1.680 ;
        RECT  1.720 2.040 2.900 2.200 ;
        RECT  2.740 1.120 2.900 2.200 ;
        RECT  2.740 1.430 3.280 1.710 ;
        RECT  1.780 1.120 2.900 1.280 ;
        RECT  1.780 0.640 1.940 1.280 ;
        RECT  1.290 2.240 1.560 2.520 ;
        RECT  1.400 0.640 1.560 2.520 ;
        RECT  1.400 1.520 2.340 1.680 ;
        RECT  1.300 0.640 1.560 0.920 ;
    END
END DELDKHD

MACRO DFCLRBEHD
    CLASS CORE ;
    FOREIGN DFCLRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.120 1.740 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.350 4.390 1.630 ;
        RECT  4.100 1.240 4.300 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.580 11.500 2.120 ;
        RECT  11.280 1.840 11.500 2.120 ;
        RECT  11.280 0.580 11.500 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 1.900 2.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 1.300 10.300 2.120 ;
        RECT  10.260 0.440 10.460 1.500 ;
        RECT  10.180 0.440 10.460 0.660 ;
        END
    END Q
    PIN LD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.820 0.700 2.640 ;
        RECT  3.100 1.500 3.260 2.640 ;
        RECT  0.500 2.480 3.260 2.640 ;
        RECT  3.100 1.500 3.420 1.780 ;
        RECT  0.480 1.820 0.700 2.100 ;
        END
    END LD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.280 4.530 0.400 ;
        RECT  7.900 -0.280 8.180 0.420 ;
        RECT  9.380 -0.280 9.660 0.420 ;
        RECT  10.760 -0.280 10.980 0.660 ;
        RECT  0.000 -0.280 11.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 2.800 2.660 3.480 ;
        RECT  4.440 2.800 4.720 3.480 ;
        RECT  7.770 2.800 8.050 3.480 ;
        RECT  8.820 2.800 9.560 3.480 ;
        RECT  10.700 2.620 10.980 3.480 ;
        RECT  0.000 2.920 11.600 3.480 ;
        RECT  0.850 2.800 1.130 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.860 2.600 6.850 2.760 ;
        RECT  6.690 2.160 6.850 2.760 ;
        RECT  3.620 2.480 3.900 2.730 ;
        RECT  9.780 2.300 10.120 2.720 ;
        RECT  8.910 2.480 10.120 2.640 ;
        RECT  5.480 2.300 6.020 2.640 ;
        RECT  3.620 2.480 6.020 2.640 ;
        RECT  8.910 1.860 9.070 2.640 ;
        RECT  9.780 2.300 11.080 2.460 ;
        RECT  10.920 1.210 11.080 2.460 ;
        RECT  6.690 2.160 7.230 2.320 ;
        RECT  7.070 1.860 7.230 2.320 ;
        RECT  9.780 0.860 9.940 2.720 ;
        RECT  5.860 0.460 6.020 2.760 ;
        RECT  7.070 1.860 9.070 2.020 ;
        RECT  9.770 0.860 10.100 1.080 ;
        RECT  5.740 0.460 6.020 0.680 ;
        RECT  9.320 0.580 9.480 2.080 ;
        RECT  9.320 1.340 9.620 1.620 ;
        RECT  8.780 0.580 9.480 0.740 ;
        RECT  6.180 2.180 6.530 2.440 ;
        RECT  6.180 0.460 6.340 2.440 ;
        RECT  8.980 1.140 9.140 1.660 ;
        RECT  6.820 1.140 9.140 1.300 ;
        RECT  6.820 0.460 6.980 1.300 ;
        RECT  6.180 0.460 6.980 0.620 ;
        RECT  8.340 0.580 8.620 0.980 ;
        RECT  7.140 0.580 8.620 0.740 ;
        RECT  7.140 0.460 7.740 0.740 ;
        RECT  7.100 2.480 7.630 2.640 ;
        RECT  8.340 2.180 8.620 2.520 ;
        RECT  7.470 2.360 8.620 2.520 ;
        RECT  6.500 1.460 6.900 1.980 ;
        RECT  6.500 1.460 8.480 1.620 ;
        RECT  6.500 0.840 6.660 1.980 ;
        RECT  1.460 2.160 2.710 2.320 ;
        RECT  2.550 0.780 2.710 2.320 ;
        RECT  3.460 2.000 3.740 2.280 ;
        RECT  3.580 0.560 3.740 2.280 ;
        RECT  5.540 0.880 5.700 2.080 ;
        RECT  5.420 0.440 5.580 1.040 ;
        RECT  1.980 0.780 3.740 0.940 ;
        RECT  3.580 0.560 4.880 0.720 ;
        RECT  4.720 0.440 5.580 0.600 ;
        RECT  5.060 0.760 5.220 2.320 ;
        RECT  5.060 1.380 5.360 1.660 ;
        RECT  3.960 2.150 4.880 2.310 ;
        RECT  4.720 0.920 4.880 2.310 ;
        RECT  3.960 0.920 4.880 1.080 ;
        RECT  1.180 0.680 1.460 0.900 ;
        RECT  1.300 0.460 1.460 0.900 ;
        RECT  1.300 0.460 3.180 0.620 ;
        RECT  0.160 0.910 0.320 2.520 ;
        RECT  2.220 1.100 2.380 1.560 ;
        RECT  0.160 1.100 2.380 1.260 ;
    END
END DFCLRBEHD

MACRO DFCLRBHHD
    CLASS CORE ;
    FOREIGN DFCLRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.120 1.740 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.350 4.390 1.630 ;
        RECT  4.100 1.240 4.300 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.100 0.840 12.300 2.360 ;
        RECT  11.960 2.080 12.300 2.360 ;
        RECT  11.960 0.840 12.300 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 1.900 2.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.960 11.100 2.260 ;
        RECT  10.840 1.980 11.100 2.260 ;
        RECT  10.840 0.960 11.100 1.240 ;
        END
    END Q
    PIN LD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.820 0.700 2.640 ;
        RECT  3.100 1.500 3.260 2.640 ;
        RECT  0.500 2.480 3.260 2.640 ;
        RECT  3.100 1.500 3.420 1.780 ;
        RECT  0.480 1.820 0.700 2.100 ;
        END
    END LD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.250 -0.280 4.530 0.400 ;
        RECT  7.900 -0.280 8.180 0.420 ;
        RECT  8.760 -0.280 9.040 0.420 ;
        RECT  10.220 -0.280 10.500 0.400 ;
        RECT  11.340 -0.280 11.620 0.400 ;
        RECT  12.420 -0.280 12.700 0.580 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 2.800 2.660 3.480 ;
        RECT  4.440 2.800 4.720 3.480 ;
        RECT  7.770 2.800 8.050 3.480 ;
        RECT  8.760 2.800 9.040 3.480 ;
        RECT  10.220 2.800 10.500 3.480 ;
        RECT  11.340 2.800 11.620 3.480 ;
        RECT  12.420 2.620 12.700 3.480 ;
        RECT  0.000 2.920 12.800 3.480 ;
        RECT  0.850 2.800 1.130 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.860 2.600 6.850 2.760 ;
        RECT  6.690 2.160 6.850 2.760 ;
        RECT  3.620 2.480 3.900 2.730 ;
        RECT  5.480 2.300 6.020 2.640 ;
        RECT  8.910 2.440 11.800 2.600 ;
        RECT  11.640 0.570 11.800 2.600 ;
        RECT  3.620 2.480 6.020 2.640 ;
        RECT  8.910 1.860 9.070 2.600 ;
        RECT  6.690 2.160 7.230 2.320 ;
        RECT  7.070 1.860 7.230 2.320 ;
        RECT  5.860 0.460 6.020 2.760 ;
        RECT  7.070 1.860 9.070 2.020 ;
        RECT  9.660 0.540 9.940 0.760 ;
        RECT  9.660 0.570 11.800 0.730 ;
        RECT  5.740 0.460 6.020 0.680 ;
        RECT  9.260 1.840 9.540 2.120 ;
        RECT  9.260 0.960 9.420 2.120 ;
        RECT  9.260 1.480 10.320 1.640 ;
        RECT  9.260 0.960 9.540 1.240 ;
        RECT  6.180 2.180 6.530 2.440 ;
        RECT  6.180 0.460 6.340 2.440 ;
        RECT  8.920 1.140 9.080 1.690 ;
        RECT  6.820 1.140 9.080 1.300 ;
        RECT  6.820 0.460 6.980 1.300 ;
        RECT  6.180 0.460 6.980 0.620 ;
        RECT  8.340 0.580 8.620 0.980 ;
        RECT  7.140 0.580 8.620 0.740 ;
        RECT  7.140 0.460 7.740 0.740 ;
        RECT  7.100 2.480 7.630 2.640 ;
        RECT  8.340 2.180 8.620 2.520 ;
        RECT  7.470 2.360 8.620 2.520 ;
        RECT  6.500 1.460 6.900 1.980 ;
        RECT  6.500 1.460 8.480 1.620 ;
        RECT  6.500 0.840 6.660 1.980 ;
        RECT  1.460 2.160 2.710 2.320 ;
        RECT  2.550 0.780 2.710 2.320 ;
        RECT  3.460 2.000 3.740 2.280 ;
        RECT  3.580 0.560 3.740 2.280 ;
        RECT  5.540 0.880 5.700 2.080 ;
        RECT  5.420 0.440 5.580 1.040 ;
        RECT  1.980 0.780 3.740 0.940 ;
        RECT  3.580 0.560 4.880 0.720 ;
        RECT  4.720 0.440 5.580 0.600 ;
        RECT  5.060 0.760 5.220 2.320 ;
        RECT  5.060 1.380 5.360 1.660 ;
        RECT  3.960 2.150 4.880 2.310 ;
        RECT  4.720 0.920 4.880 2.310 ;
        RECT  3.960 0.920 4.880 1.080 ;
        RECT  1.180 0.680 1.460 0.900 ;
        RECT  1.300 0.460 1.460 0.900 ;
        RECT  1.300 0.460 3.180 0.620 ;
        RECT  0.160 0.910 0.320 2.520 ;
        RECT  2.220 1.100 2.380 1.560 ;
        RECT  0.160 1.100 2.380 1.260 ;
    END
END DFCLRBHHD

MACRO DFCRBEHD
    CLASS CORE ;
    FOREIGN DFCRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.320 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.350 2.010 1.630 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.580 9.100 2.120 ;
        RECT  8.880 1.840 9.100 2.120 ;
        RECT  8.880 0.580 9.100 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 1.960 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.880 0.440 8.080 1.100 ;
        RECT  7.880 0.900 8.300 1.100 ;
        RECT  8.100 0.900 8.300 2.120 ;
        RECT  7.760 1.840 8.300 2.120 ;
        RECT  7.780 0.440 8.080 0.660 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.870 -0.280 2.150 0.400 ;
        RECT  5.520 -0.280 5.800 0.420 ;
        RECT  7.000 -0.280 7.280 0.420 ;
        RECT  8.300 -0.280 8.580 0.580 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 2.800 1.320 3.480 ;
        RECT  2.060 2.800 2.340 3.480 ;
        RECT  5.390 2.800 5.670 3.480 ;
        RECT  6.440 2.800 7.160 3.480 ;
        RECT  8.300 2.620 8.580 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.480 2.600 4.470 2.760 ;
        RECT  4.310 2.160 4.470 2.760 ;
        RECT  7.380 2.300 7.720 2.720 ;
        RECT  6.530 2.480 7.720 2.640 ;
        RECT  3.480 0.460 3.640 2.760 ;
        RECT  6.530 1.860 6.690 2.640 ;
        RECT  7.380 2.300 8.680 2.460 ;
        RECT  8.520 1.210 8.680 2.460 ;
        RECT  3.060 2.300 3.640 2.460 ;
        RECT  4.310 2.160 4.850 2.320 ;
        RECT  4.690 1.860 4.850 2.320 ;
        RECT  7.400 0.860 7.560 2.720 ;
        RECT  4.690 1.860 6.690 2.020 ;
        RECT  7.390 0.860 7.720 1.080 ;
        RECT  3.360 0.460 3.640 0.680 ;
        RECT  6.940 0.580 7.100 2.080 ;
        RECT  6.940 1.340 7.240 1.620 ;
        RECT  6.400 0.580 7.100 0.740 ;
        RECT  3.800 2.180 4.150 2.440 ;
        RECT  3.800 0.460 3.960 2.440 ;
        RECT  6.600 1.140 6.760 1.660 ;
        RECT  4.440 1.140 6.760 1.300 ;
        RECT  4.440 0.460 4.600 1.300 ;
        RECT  3.800 0.460 4.600 0.620 ;
        RECT  5.960 0.580 6.240 0.980 ;
        RECT  4.760 0.580 6.240 0.740 ;
        RECT  4.760 0.460 5.360 0.740 ;
        RECT  4.720 2.480 5.250 2.640 ;
        RECT  5.960 2.180 6.240 2.520 ;
        RECT  5.090 2.360 6.240 2.520 ;
        RECT  4.120 1.460 4.520 1.980 ;
        RECT  4.120 1.460 6.100 1.620 ;
        RECT  4.120 0.840 4.280 1.980 ;
        RECT  0.520 2.240 0.820 2.460 ;
        RECT  0.520 0.560 0.680 2.460 ;
        RECT  3.160 0.880 3.320 2.080 ;
        RECT  3.040 0.440 3.200 1.040 ;
        RECT  0.520 0.560 2.500 0.720 ;
        RECT  2.340 0.440 3.200 0.600 ;
        RECT  2.680 0.760 2.840 2.340 ;
        RECT  2.680 1.380 2.980 1.660 ;
        RECT  1.580 2.200 2.500 2.360 ;
        RECT  2.340 0.920 2.500 2.360 ;
        RECT  1.580 0.920 2.500 1.080 ;
    END
END DFCRBEHD

MACRO DFCRBHHD
    CLASS CORE ;
    FOREIGN DFCRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.320 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.350 2.010 1.630 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.840 9.900 2.360 ;
        RECT  9.560 2.080 9.900 2.360 ;
        RECT  9.560 0.840 9.900 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 1.960 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.960 8.700 2.260 ;
        RECT  8.440 1.980 8.700 2.260 ;
        RECT  8.440 0.960 8.700 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.870 -0.280 2.150 0.400 ;
        RECT  5.520 -0.280 5.800 0.420 ;
        RECT  6.360 -0.280 6.640 0.420 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  8.940 -0.280 9.220 0.400 ;
        RECT  10.020 -0.280 10.300 0.580 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 2.800 1.320 3.480 ;
        RECT  2.060 2.800 2.340 3.480 ;
        RECT  5.390 2.800 5.670 3.480 ;
        RECT  6.360 2.800 6.640 3.480 ;
        RECT  7.820 2.800 8.100 3.480 ;
        RECT  8.940 2.800 9.220 3.480 ;
        RECT  10.020 2.620 10.300 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.480 2.600 4.470 2.760 ;
        RECT  4.310 2.160 4.470 2.760 ;
        RECT  6.450 2.440 9.400 2.600 ;
        RECT  9.240 0.560 9.400 2.600 ;
        RECT  3.480 0.460 3.640 2.760 ;
        RECT  3.060 2.300 3.640 2.460 ;
        RECT  6.450 1.860 6.610 2.600 ;
        RECT  4.310 2.160 4.850 2.320 ;
        RECT  4.690 1.860 4.850 2.320 ;
        RECT  4.690 1.860 6.610 2.020 ;
        RECT  7.260 0.540 7.540 0.760 ;
        RECT  7.260 0.560 9.400 0.720 ;
        RECT  3.360 0.460 3.640 0.680 ;
        RECT  6.860 1.840 7.140 2.120 ;
        RECT  6.860 0.960 7.020 2.120 ;
        RECT  6.860 1.480 7.920 1.640 ;
        RECT  6.860 0.960 7.140 1.240 ;
        RECT  3.800 2.180 4.150 2.440 ;
        RECT  3.800 0.460 3.960 2.440 ;
        RECT  6.520 1.140 6.680 1.690 ;
        RECT  4.440 1.140 6.680 1.300 ;
        RECT  4.440 0.460 4.600 1.300 ;
        RECT  3.800 0.460 4.600 0.620 ;
        RECT  5.960 0.580 6.240 0.980 ;
        RECT  4.760 0.580 6.240 0.740 ;
        RECT  4.760 0.460 5.360 0.740 ;
        RECT  4.720 2.480 5.250 2.640 ;
        RECT  5.960 2.180 6.240 2.520 ;
        RECT  5.090 2.360 6.240 2.520 ;
        RECT  4.120 1.460 4.520 1.980 ;
        RECT  4.120 1.460 6.100 1.620 ;
        RECT  4.120 0.840 4.280 1.980 ;
        RECT  0.520 2.240 0.820 2.460 ;
        RECT  0.520 0.560 0.680 2.460 ;
        RECT  3.160 0.880 3.320 2.080 ;
        RECT  3.040 0.440 3.200 1.040 ;
        RECT  0.520 0.560 2.500 0.720 ;
        RECT  2.340 0.440 3.200 0.600 ;
        RECT  2.680 0.760 2.840 2.340 ;
        RECT  2.680 1.380 2.980 1.660 ;
        RECT  1.580 2.200 2.500 2.360 ;
        RECT  2.340 0.920 2.500 2.360 ;
        RECT  1.580 0.920 2.500 1.080 ;
    END
END DFCRBHHD

MACRO DFECHD
    CLASS CORE ;
    FOREIGN DFECHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 0.840 10.300 2.120 ;
        RECT  10.060 1.840 10.300 2.120 ;
        RECT  10.060 0.840 10.300 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.880 9.180 1.160 ;
        RECT  8.900 1.840 9.180 2.120 ;
        RECT  8.900 0.880 9.100 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 3.420 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  7.620 -0.280 7.900 0.420 ;
        RECT  9.480 -0.280 9.760 0.860 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 3.520 3.480 ;
        RECT  6.570 2.800 6.850 3.480 ;
        RECT  7.340 2.800 8.100 3.480 ;
        RECT  9.520 2.800 9.800 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  8.380 2.420 8.740 2.660 ;
        RECT  8.580 0.460 8.740 2.660 ;
        RECT  4.280 2.300 4.820 2.640 ;
        RECT  2.440 2.480 4.820 2.640 ;
        RECT  7.770 2.420 9.860 2.580 ;
        RECT  9.700 1.210 9.860 2.580 ;
        RECT  2.440 1.810 2.600 2.640 ;
        RECT  7.770 1.880 7.930 2.580 ;
        RECT  5.490 2.160 6.700 2.320 ;
        RECT  6.540 1.880 6.700 2.320 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  6.540 1.880 7.930 2.040 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  8.580 0.460 8.940 0.620 ;
        RECT  8.120 0.880 8.280 2.120 ;
        RECT  8.120 1.340 8.420 1.620 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.780 1.060 7.940 1.660 ;
        RECT  5.620 1.060 7.940 1.220 ;
        RECT  5.620 0.460 5.780 1.220 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  5.300 1.820 5.700 1.980 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  5.300 1.380 7.560 1.540 ;
        RECT  7.060 0.580 7.340 0.900 ;
        RECT  5.940 0.580 7.340 0.740 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  5.810 2.480 6.410 2.760 ;
        RECT  5.810 2.480 7.340 2.640 ;
        RECT  7.060 2.200 7.340 2.640 ;
        RECT  1.490 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.740 0.720 ;
        RECT  3.580 0.440 4.380 0.600 ;
        RECT  3.860 0.840 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.880 3.680 2.310 ;
        RECT  2.760 0.880 3.680 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFECHD

MACRO DFEEHD
    CLASS CORE ;
    FOREIGN DFEEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.310 3.160 1.590 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.840 10.700 2.360 ;
        RECT  10.460 2.080 10.700 2.360 ;
        RECT  10.460 0.840 10.700 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.960 9.580 1.240 ;
        RECT  9.300 1.840 9.580 2.120 ;
        RECT  9.300 0.960 9.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 3.480 0.400 ;
        RECT  6.760 -0.280 7.040 0.420 ;
        RECT  7.680 -0.280 7.960 0.420 ;
        RECT  9.020 -0.280 9.300 0.620 ;
        RECT  9.880 -0.280 10.160 0.580 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 3.580 3.480 ;
        RECT  6.630 2.800 6.910 3.480 ;
        RECT  7.500 2.800 7.780 3.480 ;
        RECT  8.410 2.800 8.690 3.480 ;
        RECT  9.880 2.620 10.160 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.720 2.600 5.710 2.760 ;
        RECT  5.550 2.160 5.710 2.760 ;
        RECT  4.340 2.300 4.880 2.640 ;
        RECT  2.440 2.480 4.880 2.640 ;
        RECT  7.830 2.420 9.460 2.580 ;
        RECT  2.440 1.810 2.600 2.640 ;
        RECT  10.100 1.210 10.260 2.440 ;
        RECT  9.300 2.280 10.260 2.440 ;
        RECT  8.660 0.460 8.820 2.580 ;
        RECT  7.830 1.880 7.990 2.580 ;
        RECT  5.550 2.160 6.760 2.320 ;
        RECT  6.600 1.880 6.760 2.320 ;
        RECT  4.720 0.460 4.880 2.760 ;
        RECT  6.600 1.880 7.990 2.040 ;
        RECT  8.500 0.460 8.820 0.680 ;
        RECT  4.600 0.460 4.880 0.680 ;
        RECT  8.180 0.880 8.340 2.120 ;
        RECT  8.180 1.340 8.480 1.620 ;
        RECT  5.040 2.180 5.390 2.440 ;
        RECT  5.040 0.460 5.200 2.440 ;
        RECT  7.840 1.060 8.000 1.660 ;
        RECT  5.680 1.060 8.000 1.220 ;
        RECT  5.680 0.460 5.840 1.220 ;
        RECT  5.040 0.460 5.840 0.620 ;
        RECT  5.360 1.820 5.760 1.980 ;
        RECT  5.360 0.840 5.520 1.980 ;
        RECT  5.360 1.380 7.620 1.540 ;
        RECT  7.120 0.580 7.400 0.900 ;
        RECT  6.000 0.580 7.400 0.740 ;
        RECT  6.000 0.460 6.600 0.740 ;
        RECT  5.870 2.480 6.470 2.760 ;
        RECT  5.870 2.480 7.400 2.640 ;
        RECT  7.120 2.200 7.400 2.640 ;
        RECT  1.490 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.400 0.880 4.560 2.080 ;
        RECT  4.280 0.440 4.440 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.800 0.720 ;
        RECT  3.640 0.440 4.440 0.600 ;
        RECT  3.920 0.840 4.080 2.320 ;
        RECT  3.920 1.380 4.220 1.660 ;
        RECT  2.820 2.150 3.740 2.310 ;
        RECT  3.580 0.880 3.740 2.310 ;
        RECT  2.820 0.880 3.740 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFEEHD

MACRO DFEHHD
    CLASS CORE ;
    FOREIGN DFEHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.310 3.160 1.590 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.840 11.100 2.360 ;
        RECT  10.760 2.080 11.100 2.360 ;
        RECT  10.760 0.840 11.100 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.960 9.900 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 3.480 0.400 ;
        RECT  6.760 -0.280 7.040 0.420 ;
        RECT  7.680 -0.280 7.960 0.420 ;
        RECT  9.140 -0.280 9.420 0.580 ;
        RECT  10.180 -0.280 10.460 0.580 ;
        RECT  11.220 -0.280 11.500 0.580 ;
        RECT  0.000 -0.280 11.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 3.580 3.480 ;
        RECT  6.630 2.800 6.910 3.480 ;
        RECT  7.640 2.800 7.920 3.480 ;
        RECT  9.140 2.620 9.420 3.480 ;
        RECT  10.180 2.620 10.460 3.480 ;
        RECT  11.220 2.620 11.500 3.480 ;
        RECT  0.000 2.920 11.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.720 2.600 5.710 2.760 ;
        RECT  5.550 2.160 5.710 2.760 ;
        RECT  4.340 2.300 4.880 2.640 ;
        RECT  2.440 2.480 4.880 2.640 ;
        RECT  7.830 2.420 8.940 2.580 ;
        RECT  8.780 0.460 8.940 2.580 ;
        RECT  2.440 1.810 2.600 2.640 ;
        RECT  10.400 1.210 10.560 2.440 ;
        RECT  8.780 2.280 10.560 2.440 ;
        RECT  7.830 1.880 7.990 2.580 ;
        RECT  5.550 2.160 6.760 2.320 ;
        RECT  6.600 1.880 6.760 2.320 ;
        RECT  4.720 0.460 4.880 2.760 ;
        RECT  6.600 1.880 7.990 2.040 ;
        RECT  8.620 0.460 8.940 0.680 ;
        RECT  4.600 0.460 4.880 0.680 ;
        RECT  8.300 0.880 8.460 2.160 ;
        RECT  8.260 1.840 8.460 2.120 ;
        RECT  8.300 1.340 8.600 1.620 ;
        RECT  5.040 2.180 5.390 2.440 ;
        RECT  5.040 0.460 5.200 2.440 ;
        RECT  7.840 1.060 8.000 1.660 ;
        RECT  5.680 1.060 8.000 1.220 ;
        RECT  5.680 0.460 5.840 1.220 ;
        RECT  5.040 0.460 5.840 0.620 ;
        RECT  5.360 1.820 5.760 1.980 ;
        RECT  5.360 0.840 5.520 1.980 ;
        RECT  5.360 1.380 7.620 1.540 ;
        RECT  7.120 0.580 7.400 0.900 ;
        RECT  6.000 0.580 7.400 0.740 ;
        RECT  6.000 0.460 6.600 0.740 ;
        RECT  5.870 2.480 6.470 2.760 ;
        RECT  5.870 2.480 7.400 2.640 ;
        RECT  7.120 2.200 7.400 2.640 ;
        RECT  1.490 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.400 0.880 4.560 2.080 ;
        RECT  4.280 0.440 4.440 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.800 0.720 ;
        RECT  3.640 0.440 4.440 0.600 ;
        RECT  3.920 0.840 4.080 2.320 ;
        RECT  3.920 1.380 4.220 1.660 ;
        RECT  2.820 2.150 3.740 2.310 ;
        RECT  3.580 0.880 3.740 2.310 ;
        RECT  2.820 0.880 3.740 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFEHHD

MACRO DFEKHD
    CLASS CORE ;
    FOREIGN DFEKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.720 0.960 12.920 1.240 ;
        RECT  11.720 1.840 12.920 2.120 ;
        RECT  12.100 0.960 12.300 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.640 0.960 10.840 1.240 ;
        RECT  9.640 1.840 10.840 2.120 ;
        RECT  10.100 0.960 10.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  6.800 -0.280 7.080 0.420 ;
        RECT  7.600 -0.280 7.880 0.420 ;
        RECT  9.060 -0.280 9.340 0.580 ;
        RECT  10.100 -0.280 10.380 0.580 ;
        RECT  11.140 -0.280 11.420 0.580 ;
        RECT  12.180 -0.280 12.460 0.580 ;
        RECT  13.220 -0.280 13.500 0.580 ;
        RECT  0.000 -0.280 13.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 3.620 3.480 ;
        RECT  6.790 2.800 7.070 3.480 ;
        RECT  7.560 2.800 7.840 3.480 ;
        RECT  9.060 2.620 9.340 3.480 ;
        RECT  10.100 2.620 10.380 3.480 ;
        RECT  11.140 2.620 11.420 3.480 ;
        RECT  12.180 2.620 12.460 3.480 ;
        RECT  13.220 2.620 13.500 3.480 ;
        RECT  0.000 2.920 13.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.760 2.600 5.750 2.760 ;
        RECT  5.590 2.160 5.750 2.760 ;
        RECT  4.380 2.300 4.920 2.640 ;
        RECT  2.410 2.480 4.920 2.640 ;
        RECT  7.750 2.420 8.860 2.580 ;
        RECT  8.700 0.460 8.860 2.580 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  11.380 1.210 11.540 2.440 ;
        RECT  8.700 2.280 11.540 2.440 ;
        RECT  7.750 1.880 7.910 2.580 ;
        RECT  5.590 2.160 6.120 2.320 ;
        RECT  5.960 1.880 6.120 2.320 ;
        RECT  4.760 0.460 4.920 2.760 ;
        RECT  5.960 1.880 7.910 2.040 ;
        RECT  8.540 0.460 8.860 0.680 ;
        RECT  4.640 0.460 4.920 0.680 ;
        RECT  8.220 0.880 8.380 2.160 ;
        RECT  8.180 1.840 8.380 2.120 ;
        RECT  8.220 1.340 8.540 1.620 ;
        RECT  5.080 2.180 5.430 2.440 ;
        RECT  5.080 0.460 5.240 2.440 ;
        RECT  7.900 1.160 8.060 1.660 ;
        RECT  5.720 1.160 8.060 1.320 ;
        RECT  5.720 0.460 5.880 1.320 ;
        RECT  5.080 0.460 5.880 0.620 ;
        RECT  5.400 1.480 5.800 1.980 ;
        RECT  5.400 1.480 7.660 1.640 ;
        RECT  5.400 0.840 5.560 1.980 ;
        RECT  7.160 0.580 7.440 0.980 ;
        RECT  6.040 0.580 7.440 0.740 ;
        RECT  6.040 0.460 6.640 0.740 ;
        RECT  5.910 2.480 6.570 2.760 ;
        RECT  6.290 2.340 6.570 2.760 ;
        RECT  7.160 2.200 7.440 2.510 ;
        RECT  6.290 2.350 7.440 2.510 ;
        RECT  1.490 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.440 0.880 4.600 2.080 ;
        RECT  4.320 0.560 4.480 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 4.480 0.720 ;
        RECT  3.960 0.880 4.120 2.320 ;
        RECT  3.960 1.380 4.260 1.660 ;
        RECT  3.940 0.880 4.160 1.160 ;
        RECT  2.740 2.150 3.780 2.310 ;
        RECT  3.620 0.880 3.780 2.310 ;
        RECT  2.740 0.880 3.780 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFEKHD

MACRO DFERBCHD
    CLASS CORE ;
    FOREIGN DFERBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.200 8.090 1.660 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.880 1.840 11.100 2.120 ;
        RECT  10.900 0.920 11.100 2.160 ;
        RECT  10.880 0.960 11.100 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.980 10.060 2.060 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.060 -0.280 3.340 0.400 ;
        RECT  6.900 -0.280 7.180 0.400 ;
        RECT  7.980 -0.280 8.260 0.400 ;
        RECT  8.820 -0.280 9.100 0.400 ;
        RECT  10.300 -0.280 10.580 0.940 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.220 2.800 3.500 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  7.500 2.800 7.780 3.480 ;
        RECT  8.620 2.800 8.900 3.480 ;
        RECT  10.260 2.620 10.540 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  4.260 2.300 4.800 2.640 ;
        RECT  2.410 2.480 4.800 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  9.380 2.220 10.630 2.380 ;
        RECT  10.470 1.290 10.630 2.380 ;
        RECT  5.710 2.160 9.540 2.320 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  9.380 0.440 9.540 2.380 ;
        RECT  10.470 1.340 10.680 1.620 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  9.380 0.440 9.700 0.600 ;
        RECT  9.060 2.600 9.400 2.760 ;
        RECT  8.020 2.480 9.220 2.640 ;
        RECT  9.060 0.880 9.220 1.760 ;
        RECT  8.800 0.880 9.220 1.160 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  8.540 1.350 8.700 1.900 ;
        RECT  6.040 1.500 7.540 1.660 ;
        RECT  7.380 0.880 7.540 1.660 ;
        RECT  8.470 0.880 8.630 1.510 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  7.380 0.880 8.630 1.040 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  6.360 1.820 8.380 1.980 ;
        RECT  6.440 0.560 7.600 0.720 ;
        RECT  7.340 0.440 7.600 0.720 ;
        RECT  5.970 0.460 6.600 0.620 ;
        RECT  6.030 2.480 7.390 2.640 ;
        RECT  6.360 0.880 7.220 1.160 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.320 0.880 4.480 2.080 ;
        RECT  4.160 0.440 4.320 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.660 0.720 ;
        RECT  3.500 0.440 4.320 0.600 ;
        RECT  3.840 0.760 4.000 2.320 ;
        RECT  3.840 1.380 4.140 1.660 ;
        RECT  2.740 2.160 3.660 2.320 ;
        RECT  3.500 0.880 3.660 2.320 ;
        RECT  2.740 0.880 3.660 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERBCHD

MACRO DFERBEHD
    CLASS CORE ;
    FOREIGN DFERBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.200 8.090 1.660 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.280 1.840 11.500 2.120 ;
        RECT  11.300 0.920 11.500 2.160 ;
        RECT  11.280 0.960 11.500 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 1.840 10.380 2.120 ;
        RECT  10.100 1.020 10.460 1.240 ;
        RECT  10.100 0.980 10.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.060 -0.280 3.340 0.400 ;
        RECT  6.900 -0.280 7.180 0.400 ;
        RECT  8.040 -0.280 8.320 0.400 ;
        RECT  9.320 -0.280 9.600 0.580 ;
        RECT  10.700 -0.280 10.980 0.580 ;
        RECT  0.000 -0.280 11.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.220 2.800 3.500 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  7.500 2.800 7.780 3.480 ;
        RECT  8.700 2.800 8.980 3.480 ;
        RECT  10.700 2.620 10.980 3.480 ;
        RECT  0.000 2.920 11.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  4.260 2.300 4.800 2.640 ;
        RECT  2.410 2.480 4.800 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  9.780 2.300 11.030 2.460 ;
        RECT  10.870 1.340 11.030 2.460 ;
        RECT  5.710 2.160 9.940 2.320 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  9.780 0.440 9.940 2.460 ;
        RECT  10.870 1.340 11.080 1.620 ;
        RECT  9.780 0.440 10.120 0.750 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  9.460 0.880 9.620 1.480 ;
        RECT  9.040 0.880 9.620 1.160 ;
        RECT  9.130 2.480 9.460 2.740 ;
        RECT  8.020 2.480 9.460 2.640 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  8.720 1.440 9.020 1.720 ;
        RECT  6.040 1.500 7.540 1.660 ;
        RECT  7.380 0.880 7.540 1.660 ;
        RECT  8.720 0.880 8.880 1.720 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  7.380 0.880 8.880 1.040 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  6.360 1.820 8.380 1.980 ;
        RECT  6.440 0.560 7.600 0.720 ;
        RECT  7.340 0.440 7.600 0.720 ;
        RECT  5.970 0.460 6.600 0.620 ;
        RECT  6.030 2.480 7.390 2.640 ;
        RECT  6.360 0.880 7.220 1.160 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.320 0.880 4.480 2.080 ;
        RECT  4.160 0.440 4.320 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.660 0.720 ;
        RECT  3.500 0.440 4.320 0.600 ;
        RECT  3.840 0.760 4.000 2.320 ;
        RECT  3.840 1.380 4.140 1.660 ;
        RECT  2.740 2.160 3.660 2.320 ;
        RECT  3.500 0.880 3.660 2.320 ;
        RECT  2.740 0.880 3.660 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERBEHD

MACRO DFERBHHD
    CLASS CORE ;
    FOREIGN DFERBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.200 8.090 1.660 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.100 0.920 12.300 2.160 ;
        RECT  11.920 1.840 12.300 2.160 ;
        RECT  11.920 0.920 12.300 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.960 11.100 2.120 ;
        RECT  10.880 1.840 11.100 2.120 ;
        RECT  10.880 0.960 11.100 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.060 -0.280 3.340 0.400 ;
        RECT  6.900 -0.280 7.180 0.400 ;
        RECT  7.980 -0.280 8.640 0.580 ;
        RECT  10.300 -0.280 10.580 0.580 ;
        RECT  11.340 -0.280 11.620 0.580 ;
        RECT  12.380 -0.280 12.660 0.580 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.220 2.800 3.500 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  7.480 2.800 7.760 3.480 ;
        RECT  8.400 2.620 8.680 3.480 ;
        RECT  9.440 2.620 9.720 3.480 ;
        RECT  10.300 2.620 10.580 3.480 ;
        RECT  11.340 2.620 11.620 3.480 ;
        RECT  12.380 2.620 12.660 3.480 ;
        RECT  0.000 2.920 12.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  4.260 2.300 4.800 2.640 ;
        RECT  2.410 2.480 4.800 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  7.570 2.300 11.670 2.460 ;
        RECT  11.510 1.340 11.670 2.460 ;
        RECT  5.710 2.160 7.730 2.320 ;
        RECT  9.840 2.020 10.120 2.460 ;
        RECT  9.960 0.780 10.120 2.460 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  11.510 1.340 11.720 1.620 ;
        RECT  9.840 0.780 10.120 1.060 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  8.880 1.950 9.680 2.110 ;
        RECT  9.520 0.490 9.680 2.110 ;
        RECT  9.520 1.460 9.800 1.740 ;
        RECT  9.200 0.490 9.680 0.650 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  9.160 0.880 9.320 1.670 ;
        RECT  6.040 1.500 7.540 1.660 ;
        RECT  7.380 0.880 7.540 1.660 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  7.380 0.880 9.320 1.040 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  8.060 1.820 8.340 2.140 ;
        RECT  6.360 1.820 8.340 1.980 ;
        RECT  6.440 0.560 7.600 0.720 ;
        RECT  7.340 0.440 7.600 0.720 ;
        RECT  5.970 0.460 6.600 0.620 ;
        RECT  6.030 2.480 7.390 2.640 ;
        RECT  6.360 0.880 7.220 1.160 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.320 0.880 4.480 2.080 ;
        RECT  4.160 0.440 4.320 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.660 0.720 ;
        RECT  3.500 0.440 4.320 0.600 ;
        RECT  3.840 0.760 4.000 2.320 ;
        RECT  3.840 1.380 4.140 1.660 ;
        RECT  2.740 2.160 3.660 2.320 ;
        RECT  3.500 0.880 3.660 2.320 ;
        RECT  2.740 0.880 3.660 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERBHHD

MACRO DFERBKHD
    CLASS CORE ;
    FOREIGN DFERBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.200 8.700 1.960 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.200 3.100 1.800 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.920 0.960 14.120 1.240 ;
        RECT  12.920 1.840 14.120 2.120 ;
        RECT  13.300 0.960 13.500 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.840 0.960 12.040 1.240 ;
        RECT  10.840 1.840 12.040 2.120 ;
        RECT  11.300 0.960 11.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  7.570 -0.280 8.170 0.460 ;
        RECT  8.390 -0.280 8.670 0.580 ;
        RECT  10.260 -0.280 10.540 0.580 ;
        RECT  11.300 -0.280 11.580 0.580 ;
        RECT  12.340 -0.280 12.620 0.580 ;
        RECT  13.380 -0.280 13.660 0.580 ;
        RECT  14.420 -0.280 14.700 0.580 ;
        RECT  0.000 -0.280 14.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.340 2.800 3.620 3.480 ;
        RECT  6.460 2.800 6.740 3.480 ;
        RECT  7.560 2.800 7.840 3.480 ;
        RECT  8.320 2.800 8.600 3.480 ;
        RECT  9.400 2.620 9.680 3.480 ;
        RECT  10.260 2.620 10.540 3.480 ;
        RECT  11.300 2.620 11.580 3.480 ;
        RECT  12.340 2.620 12.620 3.480 ;
        RECT  13.380 2.620 13.660 3.480 ;
        RECT  14.420 2.620 14.700 3.480 ;
        RECT  0.000 2.920 14.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.760 2.600 5.730 2.760 ;
        RECT  5.570 2.160 5.730 2.760 ;
        RECT  4.380 2.300 4.920 2.640 ;
        RECT  2.410 2.480 4.920 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  7.690 2.300 12.670 2.460 ;
        RECT  12.510 1.340 12.670 2.460 ;
        RECT  5.570 2.160 7.850 2.320 ;
        RECT  9.800 2.020 10.080 2.460 ;
        RECT  9.920 0.960 10.080 2.460 ;
        RECT  4.760 0.460 4.920 2.760 ;
        RECT  12.510 1.340 12.720 1.620 ;
        RECT  9.800 0.960 10.080 1.240 ;
        RECT  4.600 0.460 4.920 0.680 ;
        RECT  8.880 1.950 9.640 2.110 ;
        RECT  9.480 0.490 9.640 2.110 ;
        RECT  8.880 1.890 9.160 2.110 ;
        RECT  9.480 1.460 9.760 1.740 ;
        RECT  9.190 0.490 9.640 0.650 ;
        RECT  5.080 2.220 5.410 2.440 ;
        RECT  5.080 0.440 5.240 2.440 ;
        RECT  9.110 0.810 9.270 1.670 ;
        RECT  7.940 0.810 9.270 0.970 ;
        RECT  7.940 0.620 8.100 0.970 ;
        RECT  7.250 0.620 8.100 0.780 ;
        RECT  7.250 0.440 7.410 0.780 ;
        RECT  5.080 0.440 7.410 0.600 ;
        RECT  8.020 1.820 8.300 2.140 ;
        RECT  5.980 1.820 8.300 1.980 ;
        RECT  6.610 1.380 7.640 1.540 ;
        RECT  7.480 0.940 7.640 1.540 ;
        RECT  6.610 1.120 6.770 1.540 ;
        RECT  5.860 1.120 6.770 1.280 ;
        RECT  7.480 0.940 7.760 1.160 ;
        RECT  5.860 0.940 6.140 1.280 ;
        RECT  5.900 2.480 6.180 2.700 ;
        RECT  5.900 2.480 7.500 2.640 ;
        RECT  6.930 0.940 7.260 1.220 ;
        RECT  6.930 0.760 7.090 1.220 ;
        RECT  6.300 0.760 7.090 0.920 ;
        RECT  5.400 1.440 5.780 1.980 ;
        RECT  6.170 1.440 6.450 1.660 ;
        RECT  5.400 1.440 6.450 1.600 ;
        RECT  5.400 0.840 5.560 1.980 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.440 0.880 4.600 2.080 ;
        RECT  4.280 0.560 4.440 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 4.440 0.720 ;
        RECT  3.960 0.880 4.120 2.320 ;
        RECT  3.960 1.380 4.260 1.660 ;
        RECT  3.900 0.880 4.120 1.160 ;
        RECT  2.740 2.160 3.740 2.320 ;
        RECT  3.580 0.880 3.740 2.320 ;
        RECT  3.580 1.460 3.780 1.740 ;
        RECT  2.740 0.880 3.740 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERBKHD

MACRO DFERSBCHD
    CLASS CORE ;
    FOREIGN DFERSBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.290 0.840 8.700 1.340 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.080 1.840 12.300 2.120 ;
        RECT  12.100 0.920 12.300 2.160 ;
        RECT  12.080 0.960 12.300 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.840 11.120 2.120 ;
        RECT  10.900 1.020 11.260 1.240 ;
        RECT  10.900 0.980 11.100 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 1.380 9.900 1.960 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.060 -0.280 3.340 0.400 ;
        RECT  7.180 -0.280 7.460 0.620 ;
        RECT  8.580 -0.280 8.860 0.620 ;
        RECT  9.800 -0.280 10.080 0.620 ;
        RECT  11.500 -0.280 11.780 0.940 ;
        RECT  0.000 -0.280 12.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.220 2.800 3.500 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  8.160 2.800 8.440 3.480 ;
        RECT  9.400 2.800 9.680 3.480 ;
        RECT  10.420 2.800 10.700 3.480 ;
        RECT  11.460 2.620 11.740 3.480 ;
        RECT  0.000 2.920 12.400 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  4.260 2.300 4.800 2.640 ;
        RECT  2.410 2.480 4.800 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  10.580 2.300 11.830 2.460 ;
        RECT  11.670 1.340 11.830 2.460 ;
        RECT  5.710 2.160 10.740 2.320 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  10.580 0.440 10.740 2.460 ;
        RECT  11.670 1.340 11.880 1.620 ;
        RECT  10.580 0.440 10.920 0.750 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  10.260 0.940 10.420 1.480 ;
        RECT  9.420 0.940 10.420 1.100 ;
        RECT  9.930 2.480 10.260 2.740 ;
        RECT  8.760 2.480 10.260 2.640 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  9.200 1.500 9.360 1.920 ;
        RECT  6.040 1.500 9.360 1.660 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  6.360 1.820 9.040 1.980 ;
        RECT  6.030 2.480 7.980 2.640 ;
        RECT  6.470 1.180 7.920 1.340 ;
        RECT  7.760 0.700 7.920 1.340 ;
        RECT  6.470 0.880 6.630 1.340 ;
        RECT  6.360 0.880 6.630 1.160 ;
        RECT  6.790 0.780 7.600 1.000 ;
        RECT  6.790 0.460 6.950 1.000 ;
        RECT  5.970 0.460 6.950 0.620 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.320 0.880 4.480 2.080 ;
        RECT  4.160 0.440 4.320 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.660 0.720 ;
        RECT  3.500 0.440 4.320 0.600 ;
        RECT  3.840 0.760 4.000 2.320 ;
        RECT  3.840 1.380 4.140 1.660 ;
        RECT  2.740 2.150 3.660 2.310 ;
        RECT  3.500 0.910 3.660 2.310 ;
        RECT  2.740 0.910 3.660 1.070 ;
        RECT  2.780 0.880 3.060 1.070 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERSBCHD

MACRO DFERSBEHD
    CLASS CORE ;
    FOREIGN DFERSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.290 0.840 8.700 1.340 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.080 1.840 12.300 2.120 ;
        RECT  12.100 0.920 12.300 2.160 ;
        RECT  12.080 0.960 12.300 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.840 11.180 2.120 ;
        RECT  10.900 1.020 11.260 1.240 ;
        RECT  10.900 0.980 11.100 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 1.380 9.900 1.960 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.060 -0.280 3.340 0.400 ;
        RECT  7.180 -0.280 7.460 0.620 ;
        RECT  8.580 -0.280 8.860 0.620 ;
        RECT  9.800 -0.280 10.080 0.620 ;
        RECT  11.500 -0.280 11.780 0.580 ;
        RECT  0.000 -0.280 12.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.220 2.800 3.500 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  8.160 2.800 8.440 3.480 ;
        RECT  9.400 2.800 9.680 3.480 ;
        RECT  10.420 2.800 10.700 3.480 ;
        RECT  11.500 2.620 11.780 3.480 ;
        RECT  0.000 2.920 12.400 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  4.260 2.300 4.800 2.640 ;
        RECT  2.410 2.480 4.800 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  10.580 2.300 11.830 2.460 ;
        RECT  11.670 1.340 11.830 2.460 ;
        RECT  5.710 2.160 10.740 2.320 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  10.580 0.440 10.740 2.460 ;
        RECT  11.670 1.340 11.880 1.620 ;
        RECT  10.580 0.440 10.920 0.750 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  10.260 0.940 10.420 1.480 ;
        RECT  9.420 0.940 10.420 1.100 ;
        RECT  9.930 2.480 10.260 2.740 ;
        RECT  8.760 2.480 10.260 2.640 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  9.200 1.500 9.360 1.920 ;
        RECT  6.040 1.500 9.360 1.660 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  6.360 1.820 9.040 1.980 ;
        RECT  6.030 2.480 7.980 2.640 ;
        RECT  6.470 1.180 7.920 1.340 ;
        RECT  7.760 0.700 7.920 1.340 ;
        RECT  6.470 0.880 6.630 1.340 ;
        RECT  6.360 0.880 6.630 1.160 ;
        RECT  6.790 0.780 7.600 1.000 ;
        RECT  6.790 0.460 6.950 1.000 ;
        RECT  5.970 0.460 6.950 0.620 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.320 0.880 4.480 2.080 ;
        RECT  4.160 0.440 4.320 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.660 0.720 ;
        RECT  3.500 0.440 4.320 0.600 ;
        RECT  3.840 0.760 4.000 2.320 ;
        RECT  3.840 1.380 4.140 1.660 ;
        RECT  2.740 2.160 3.660 2.320 ;
        RECT  3.500 0.880 3.660 2.320 ;
        RECT  2.740 0.880 3.660 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERSBEHD

MACRO DFERSBHHD
    CLASS CORE ;
    FOREIGN DFERSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.620 9.120 1.900 ;
        RECT  8.900 1.440 9.100 1.940 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 0.920 13.500 2.160 ;
        RECT  13.160 1.840 13.500 2.160 ;
        RECT  13.160 0.920 13.500 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.060 0.960 12.340 1.240 ;
        RECT  12.060 1.840 12.340 2.120 ;
        RECT  12.100 0.960 12.300 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.420 10.700 1.960 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.060 -0.280 3.340 0.400 ;
        RECT  7.230 -0.280 7.450 0.680 ;
        RECT  9.000 -0.280 9.280 0.620 ;
        RECT  10.320 -0.280 10.600 0.620 ;
        RECT  11.500 -0.280 11.780 0.400 ;
        RECT  12.580 -0.280 12.860 0.580 ;
        RECT  13.620 -0.280 13.900 0.580 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.220 2.800 3.500 3.480 ;
        RECT  6.680 2.800 6.960 3.480 ;
        RECT  8.300 2.800 8.580 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  10.380 2.800 10.660 3.480 ;
        RECT  11.500 2.800 11.780 3.480 ;
        RECT  12.580 2.620 12.860 3.480 ;
        RECT  13.620 2.620 13.900 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.640 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  8.210 2.480 12.350 2.640 ;
        RECT  12.190 2.280 12.350 2.640 ;
        RECT  4.260 2.300 4.800 2.640 ;
        RECT  2.410 2.480 4.800 2.640 ;
        RECT  11.720 0.900 11.880 2.640 ;
        RECT  8.210 2.160 8.370 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  12.190 2.280 13.000 2.440 ;
        RECT  12.840 1.300 13.000 2.440 ;
        RECT  5.710 2.160 8.370 2.320 ;
        RECT  4.640 0.460 4.800 2.760 ;
        RECT  11.220 0.900 11.880 1.060 ;
        RECT  11.220 0.750 11.440 1.060 ;
        RECT  4.480 0.460 4.800 0.680 ;
        RECT  9.740 2.160 11.480 2.320 ;
        RECT  11.320 1.240 11.480 2.320 ;
        RECT  10.880 1.240 11.480 1.400 ;
        RECT  10.880 0.780 11.040 1.400 ;
        RECT  9.840 0.780 10.160 1.040 ;
        RECT  9.840 0.780 11.040 0.940 ;
        RECT  5.270 2.280 5.550 2.440 ;
        RECT  5.310 1.840 5.470 2.440 ;
        RECT  5.310 1.840 6.200 2.000 ;
        RECT  6.040 1.060 6.200 2.000 ;
        RECT  10.060 1.200 10.220 1.940 ;
        RECT  6.040 1.500 8.720 1.660 ;
        RECT  8.560 0.880 8.720 1.660 ;
        RECT  9.480 1.200 10.220 1.360 ;
        RECT  5.620 1.060 6.200 1.220 ;
        RECT  9.480 0.880 9.640 1.360 ;
        RECT  5.620 0.600 5.780 1.220 ;
        RECT  8.560 0.880 9.640 1.040 ;
        RECT  5.000 0.600 5.780 0.760 ;
        RECT  5.000 0.460 5.340 0.760 ;
        RECT  8.530 2.160 9.150 2.320 ;
        RECT  8.530 1.820 8.690 2.320 ;
        RECT  6.360 1.820 8.690 1.980 ;
        RECT  6.790 0.840 7.860 1.000 ;
        RECT  7.700 0.560 7.860 1.000 ;
        RECT  6.790 0.460 6.950 1.000 ;
        RECT  7.700 0.560 8.580 0.720 ;
        RECT  5.970 0.460 6.950 0.620 ;
        RECT  6.470 1.180 8.400 1.340 ;
        RECT  8.150 0.880 8.400 1.340 ;
        RECT  6.470 0.880 6.630 1.340 ;
        RECT  6.360 0.880 6.630 1.160 ;
        RECT  6.030 2.480 8.050 2.640 ;
        RECT  4.960 0.940 5.120 2.080 ;
        RECT  4.960 1.380 5.880 1.660 ;
        RECT  4.960 0.940 5.320 1.100 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.320 0.880 4.480 2.040 ;
        RECT  4.160 0.440 4.320 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 3.660 0.720 ;
        RECT  3.500 0.440 4.320 0.600 ;
        RECT  3.840 0.760 4.000 2.320 ;
        RECT  3.840 1.380 4.140 1.660 ;
        RECT  2.740 2.160 3.660 2.320 ;
        RECT  3.500 0.880 3.660 2.320 ;
        RECT  2.740 0.880 3.660 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERSBHHD

MACRO DFERSBKHD
    CLASS CORE ;
    FOREIGN DFERSBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.350 9.100 1.940 ;
        RECT  8.880 1.620 9.100 1.900 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.250 0.700 1.970 ;
        RECT  0.480 1.660 0.700 1.940 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.170 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.120 0.960 15.320 1.240 ;
        RECT  14.120 1.840 15.320 2.120 ;
        RECT  14.450 0.960 14.750 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.380 1.580 1.660 ;
        RECT  1.300 1.340 1.500 2.010 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.040 0.960 13.240 1.240 ;
        RECT  12.040 1.840 13.240 2.120 ;
        RECT  12.450 0.960 12.750 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.260 10.700 1.960 ;
        RECT  10.480 1.420 10.700 1.700 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 -0.280 2.700 0.400 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  7.260 -0.280 7.540 0.400 ;
        RECT  8.920 -0.280 9.200 0.620 ;
        RECT  10.240 -0.280 10.520 0.620 ;
        RECT  11.420 -0.280 11.700 0.400 ;
        RECT  12.500 -0.280 12.780 0.580 ;
        RECT  13.540 -0.280 13.820 0.580 ;
        RECT  14.580 -0.280 14.860 0.580 ;
        RECT  15.620 -0.280 15.900 0.580 ;
        RECT  0.000 -0.280 16.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.800 2.700 3.480 ;
        RECT  3.340 2.800 3.620 3.480 ;
        RECT  6.630 2.800 6.910 3.480 ;
        RECT  8.220 2.800 8.500 3.480 ;
        RECT  9.100 2.800 9.380 3.480 ;
        RECT  10.300 2.800 10.580 3.480 ;
        RECT  11.420 2.800 11.700 3.480 ;
        RECT  12.500 2.620 12.780 3.480 ;
        RECT  13.540 2.620 13.820 3.480 ;
        RECT  14.580 2.620 14.860 3.480 ;
        RECT  15.620 2.620 15.900 3.480 ;
        RECT  0.000 2.920 16.000 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.760 2.600 5.730 2.760 ;
        RECT  5.570 2.160 5.730 2.760 ;
        RECT  8.130 2.480 12.270 2.640 ;
        RECT  12.110 2.280 12.270 2.640 ;
        RECT  4.380 2.300 4.920 2.640 ;
        RECT  2.410 2.480 4.920 2.640 ;
        RECT  11.640 0.900 11.800 2.640 ;
        RECT  8.130 2.160 8.290 2.640 ;
        RECT  2.410 1.810 2.570 2.640 ;
        RECT  12.110 2.280 13.960 2.440 ;
        RECT  13.800 1.300 13.960 2.440 ;
        RECT  5.570 2.160 8.290 2.320 ;
        RECT  4.760 0.460 4.920 2.760 ;
        RECT  11.180 0.900 11.800 1.060 ;
        RECT  11.180 0.750 11.400 1.060 ;
        RECT  4.600 0.460 4.920 0.680 ;
        RECT  9.660 2.160 11.440 2.320 ;
        RECT  11.280 1.240 11.440 2.320 ;
        RECT  10.860 1.240 11.440 1.400 ;
        RECT  10.860 0.780 11.020 1.400 ;
        RECT  9.760 0.780 10.080 1.040 ;
        RECT  9.760 0.780 11.020 0.940 ;
        RECT  5.080 2.280 5.410 2.440 ;
        RECT  5.080 0.440 5.240 2.440 ;
        RECT  9.980 1.200 10.140 1.940 ;
        RECT  9.400 1.200 10.140 1.360 ;
        RECT  9.400 0.790 9.560 1.360 ;
        RECT  8.560 0.790 9.560 0.950 ;
        RECT  8.560 0.560 8.720 0.950 ;
        RECT  6.870 0.560 8.720 0.720 ;
        RECT  5.080 0.440 7.030 0.600 ;
        RECT  8.450 2.160 9.070 2.320 ;
        RECT  8.450 1.840 8.610 2.320 ;
        RECT  5.980 1.840 8.610 2.000 ;
        RECT  6.980 1.500 8.260 1.660 ;
        RECT  8.100 0.880 8.260 1.660 ;
        RECT  6.980 1.200 7.140 1.660 ;
        RECT  5.920 1.200 7.140 1.360 ;
        RECT  5.920 0.830 6.080 1.360 ;
        RECT  8.100 0.880 8.320 1.160 ;
        RECT  5.980 2.480 7.970 2.640 ;
        RECT  7.360 1.160 7.740 1.320 ;
        RECT  7.360 0.880 7.520 1.320 ;
        RECT  6.340 0.880 7.520 1.040 ;
        RECT  6.340 0.760 6.620 1.040 ;
        RECT  5.400 1.520 5.780 1.980 ;
        RECT  5.400 1.520 6.770 1.680 ;
        RECT  5.400 0.840 5.560 1.980 ;
        RECT  1.500 2.520 2.220 2.680 ;
        RECT  2.060 0.560 2.220 2.680 ;
        RECT  4.440 0.880 4.600 2.040 ;
        RECT  4.280 0.560 4.440 1.040 ;
        RECT  1.500 0.740 2.220 0.900 ;
        RECT  2.060 0.560 4.440 0.720 ;
        RECT  3.960 0.880 4.120 2.320 ;
        RECT  3.960 1.380 4.260 1.660 ;
        RECT  3.900 0.880 4.120 1.160 ;
        RECT  2.740 2.160 3.730 2.320 ;
        RECT  3.570 0.880 3.730 2.320 ;
        RECT  2.740 0.880 3.730 1.040 ;
        RECT  0.160 0.780 0.320 2.580 ;
        RECT  0.160 2.200 1.900 2.360 ;
        RECT  1.740 1.820 1.900 2.360 ;
        RECT  0.860 1.190 1.140 1.450 ;
        RECT  0.860 0.780 1.020 1.450 ;
        RECT  0.160 0.780 1.020 0.940 ;
    END
END DFERSBKHD

MACRO DFFCHD
    CLASS CORE ;
    FOREIGN DFFCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.580 8.700 2.120 ;
        RECT  8.480 1.840 8.700 2.120 ;
        RECT  8.480 0.580 8.700 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.440 7.660 0.660 ;
        RECT  7.300 0.440 7.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 -0.280 1.690 0.400 ;
        RECT  4.970 -0.280 5.250 0.420 ;
        RECT  6.450 -0.280 6.730 0.420 ;
        RECT  7.960 -0.280 8.180 0.660 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.510 2.800 1.790 3.480 ;
        RECT  4.840 2.800 5.120 3.480 ;
        RECT  5.890 2.800 6.630 3.480 ;
        RECT  7.940 2.800 8.220 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.930 2.600 3.920 2.760 ;
        RECT  3.760 2.160 3.920 2.760 ;
        RECT  6.850 2.480 7.190 2.720 ;
        RECT  5.980 2.480 8.280 2.640 ;
        RECT  8.120 1.210 8.280 2.640 ;
        RECT  2.930 0.460 3.090 2.760 ;
        RECT  6.850 0.860 7.010 2.720 ;
        RECT  5.980 1.860 6.140 2.640 ;
        RECT  2.510 2.300 3.090 2.460 ;
        RECT  3.760 2.160 4.300 2.320 ;
        RECT  4.140 1.860 4.300 2.320 ;
        RECT  4.140 1.860 6.140 2.020 ;
        RECT  6.850 0.860 7.110 1.140 ;
        RECT  2.810 0.460 3.090 0.680 ;
        RECT  6.390 0.580 6.550 2.120 ;
        RECT  6.390 1.340 6.690 1.620 ;
        RECT  5.850 0.580 6.550 0.740 ;
        RECT  3.250 2.180 3.600 2.440 ;
        RECT  3.250 0.460 3.410 2.440 ;
        RECT  6.050 1.140 6.210 1.660 ;
        RECT  3.890 1.140 6.210 1.300 ;
        RECT  3.890 0.460 4.050 1.300 ;
        RECT  3.250 0.460 4.050 0.620 ;
        RECT  5.410 0.580 5.690 0.980 ;
        RECT  4.210 0.580 5.690 0.740 ;
        RECT  4.210 0.460 4.810 0.740 ;
        RECT  4.170 2.480 4.700 2.640 ;
        RECT  5.410 2.180 5.690 2.520 ;
        RECT  4.540 2.360 5.690 2.520 ;
        RECT  3.570 1.460 3.970 1.980 ;
        RECT  3.570 1.460 5.550 1.620 ;
        RECT  3.570 0.840 3.730 1.980 ;
        RECT  0.600 0.560 0.760 2.300 ;
        RECT  2.610 0.880 2.770 2.080 ;
        RECT  2.490 0.440 2.650 1.040 ;
        RECT  0.600 0.560 2.010 0.720 ;
        RECT  1.850 0.440 2.650 0.600 ;
        RECT  2.130 0.840 2.290 2.320 ;
        RECT  2.130 1.380 2.430 1.660 ;
        RECT  1.030 2.150 1.950 2.310 ;
        RECT  1.790 0.900 1.950 2.310 ;
        RECT  1.030 0.900 1.950 1.060 ;
    END
END DFFCHD

MACRO DFFEHD
    CLASS CORE ;
    FOREIGN DFFEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.580 8.700 2.120 ;
        RECT  8.480 1.840 8.700 2.120 ;
        RECT  8.480 0.580 8.700 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.440 7.660 0.660 ;
        RECT  7.300 0.440 7.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 -0.280 1.690 0.400 ;
        RECT  4.970 -0.280 5.250 0.420 ;
        RECT  6.450 -0.280 6.730 0.420 ;
        RECT  7.900 -0.280 8.180 0.600 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.510 2.800 1.790 3.480 ;
        RECT  4.840 2.800 5.120 3.480 ;
        RECT  5.890 2.800 6.630 3.480 ;
        RECT  7.900 2.620 8.180 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.930 2.600 3.920 2.760 ;
        RECT  3.760 2.160 3.920 2.760 ;
        RECT  6.850 2.290 7.270 2.720 ;
        RECT  5.980 2.480 7.270 2.640 ;
        RECT  2.930 0.460 3.090 2.760 ;
        RECT  5.980 1.860 6.140 2.640 ;
        RECT  2.510 2.300 3.090 2.460 ;
        RECT  6.850 2.290 8.280 2.450 ;
        RECT  8.120 1.210 8.280 2.450 ;
        RECT  3.760 2.160 4.300 2.320 ;
        RECT  4.140 1.860 4.300 2.320 ;
        RECT  6.850 0.860 7.010 2.720 ;
        RECT  4.140 1.860 6.140 2.020 ;
        RECT  6.850 0.860 7.110 1.140 ;
        RECT  2.810 0.460 3.090 0.680 ;
        RECT  6.390 0.580 6.550 2.120 ;
        RECT  6.390 1.340 6.690 1.620 ;
        RECT  5.850 0.580 6.550 0.740 ;
        RECT  3.250 2.180 3.600 2.440 ;
        RECT  3.250 0.460 3.410 2.440 ;
        RECT  6.050 1.140 6.210 1.660 ;
        RECT  3.890 1.140 6.210 1.300 ;
        RECT  3.890 0.460 4.050 1.300 ;
        RECT  3.250 0.460 4.050 0.620 ;
        RECT  5.410 0.580 5.690 0.980 ;
        RECT  4.210 0.580 5.690 0.740 ;
        RECT  4.210 0.460 4.810 0.740 ;
        RECT  4.170 2.480 4.700 2.640 ;
        RECT  5.410 2.180 5.690 2.520 ;
        RECT  4.540 2.360 5.690 2.520 ;
        RECT  3.570 1.460 3.970 1.980 ;
        RECT  3.570 1.460 5.550 1.620 ;
        RECT  3.570 0.840 3.730 1.980 ;
        RECT  0.600 0.560 0.760 2.300 ;
        RECT  2.610 0.880 2.770 2.080 ;
        RECT  2.490 0.440 2.650 1.040 ;
        RECT  0.600 0.560 2.010 0.720 ;
        RECT  1.850 0.440 2.650 0.600 ;
        RECT  2.130 0.840 2.290 2.320 ;
        RECT  2.130 1.380 2.430 1.660 ;
        RECT  1.030 2.150 1.950 2.310 ;
        RECT  1.790 0.900 1.950 2.310 ;
        RECT  1.030 0.900 1.950 1.060 ;
    END
END DFFEHD

MACRO DFFHHD
    CLASS CORE ;
    FOREIGN DFFHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.350 1.590 1.630 ;
        RECT  1.300 1.240 1.500 1.780 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.960 7.500 2.120 ;
        RECT  7.120 1.840 7.500 2.120 ;
        RECT  7.120 0.960 7.500 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.880 8.700 2.120 ;
        RECT  8.240 1.840 8.700 2.120 ;
        RECT  8.240 0.880 8.700 1.160 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.450 -0.280 1.730 0.400 ;
        RECT  5.100 -0.280 5.380 0.420 ;
        RECT  6.500 -0.280 6.780 0.400 ;
        RECT  7.620 -0.280 7.900 0.400 ;
        RECT  8.700 -0.280 8.980 0.580 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.640 2.800 1.920 3.480 ;
        RECT  4.970 2.800 5.250 3.480 ;
        RECT  6.540 2.620 6.820 3.480 ;
        RECT  7.620 2.800 7.900 3.480 ;
        RECT  8.700 2.620 8.980 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.060 2.600 4.050 2.760 ;
        RECT  3.890 2.160 4.050 2.760 ;
        RECT  3.060 0.460 3.220 2.760 ;
        RECT  6.100 2.300 9.440 2.460 ;
        RECT  9.280 0.500 9.440 2.460 ;
        RECT  2.640 2.300 3.220 2.460 ;
        RECT  5.700 2.220 6.260 2.380 ;
        RECT  3.890 2.160 4.430 2.320 ;
        RECT  6.800 1.370 6.960 2.460 ;
        RECT  5.700 2.030 5.860 2.380 ;
        RECT  4.270 2.030 5.860 2.190 ;
        RECT  2.940 0.460 3.220 0.680 ;
        RECT  6.020 1.840 6.460 2.060 ;
        RECT  6.300 0.640 6.460 2.060 ;
        RECT  7.920 0.640 8.080 1.710 ;
        RECT  6.180 0.440 6.340 0.970 ;
        RECT  6.180 0.640 8.080 0.800 ;
        RECT  5.900 0.440 6.340 0.600 ;
        RECT  3.380 2.180 3.730 2.440 ;
        RECT  3.380 0.460 3.540 2.440 ;
        RECT  5.880 1.350 6.100 1.630 ;
        RECT  4.020 1.350 6.100 1.510 ;
        RECT  4.020 0.460 4.180 1.510 ;
        RECT  3.380 0.460 4.180 0.620 ;
        RECT  4.780 0.940 5.860 1.100 ;
        RECT  4.780 0.460 4.940 1.100 ;
        RECT  4.340 0.460 4.940 0.740 ;
        RECT  5.380 2.540 5.860 2.700 ;
        RECT  4.300 2.480 4.830 2.640 ;
        RECT  5.380 2.360 5.540 2.700 ;
        RECT  4.670 2.360 5.540 2.520 ;
        RECT  3.700 1.680 4.100 1.980 ;
        RECT  3.700 1.680 5.680 1.840 ;
        RECT  3.700 0.840 3.860 1.980 ;
        RECT  0.600 0.560 0.760 2.310 ;
        RECT  2.740 0.880 2.900 2.080 ;
        RECT  2.620 0.440 2.780 1.040 ;
        RECT  0.600 0.560 2.080 0.720 ;
        RECT  1.920 0.440 2.780 0.600 ;
        RECT  2.260 0.760 2.420 2.320 ;
        RECT  2.260 1.380 2.560 1.660 ;
        RECT  1.160 2.150 2.080 2.310 ;
        RECT  1.920 0.920 2.080 2.310 ;
        RECT  1.160 0.920 2.080 1.080 ;
    END
END DFFHHD

MACRO DFFKHD
    CLASS CORE ;
    FOREIGN DFFKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        RECT  1.660 1.350 1.900 1.630 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.360 0.960 8.640 1.240 ;
        RECT  7.520 1.840 8.720 2.120 ;
        RECT  8.100 0.960 8.300 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.600 0.880 10.800 1.160 ;
        RECT  9.600 1.840 10.800 2.120 ;
        RECT  10.100 0.880 10.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.280 2.120 0.400 ;
        RECT  5.300 -0.280 5.580 0.420 ;
        RECT  6.740 -0.280 7.020 0.400 ;
        RECT  7.860 -0.280 8.140 0.400 ;
        RECT  8.980 -0.280 9.260 0.400 ;
        RECT  10.060 -0.280 10.340 0.580 ;
        RECT  11.100 -0.280 11.380 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 2.800 2.120 3.480 ;
        RECT  5.400 2.800 5.680 3.480 ;
        RECT  6.940 2.620 7.220 3.480 ;
        RECT  7.980 2.620 8.260 3.480 ;
        RECT  9.020 2.620 9.300 3.480 ;
        RECT  10.060 2.620 10.340 3.480 ;
        RECT  11.100 2.620 11.380 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.260 2.600 4.250 2.760 ;
        RECT  4.090 2.160 4.250 2.760 ;
        RECT  3.260 0.460 3.420 2.760 ;
        RECT  7.180 2.300 11.840 2.460 ;
        RECT  11.680 0.500 11.840 2.460 ;
        RECT  2.840 2.300 3.420 2.460 ;
        RECT  6.160 2.280 7.340 2.440 ;
        RECT  4.090 2.160 4.630 2.320 ;
        RECT  7.180 1.400 7.340 2.460 ;
        RECT  6.160 2.000 6.320 2.440 ;
        RECT  4.470 2.000 6.320 2.160 ;
        RECT  3.140 0.460 3.420 0.680 ;
        RECT  6.480 1.840 6.680 2.120 ;
        RECT  6.520 0.640 6.680 2.120 ;
        RECT  9.280 0.640 9.440 1.710 ;
        RECT  6.360 0.640 6.680 0.870 ;
        RECT  6.360 0.640 9.440 0.800 ;
        RECT  6.180 0.440 6.580 0.660 ;
        RECT  3.580 2.180 3.930 2.440 ;
        RECT  3.580 0.460 3.740 2.440 ;
        RECT  6.080 1.260 6.360 1.580 ;
        RECT  4.220 1.260 6.360 1.420 ;
        RECT  4.220 0.460 4.380 1.420 ;
        RECT  3.580 0.460 4.380 0.620 ;
        RECT  5.840 2.600 6.320 2.760 ;
        RECT  4.500 2.480 5.030 2.640 ;
        RECT  5.840 2.340 6.000 2.760 ;
        RECT  4.870 2.340 6.000 2.500 ;
        RECT  4.980 0.940 6.060 1.100 ;
        RECT  4.980 0.460 5.140 1.100 ;
        RECT  4.540 0.460 5.140 0.740 ;
        RECT  3.900 1.580 4.300 1.980 ;
        RECT  3.900 1.580 5.880 1.740 ;
        RECT  3.900 0.840 4.060 1.980 ;
        RECT  0.600 0.560 0.760 2.300 ;
        RECT  2.940 0.880 3.100 2.080 ;
        RECT  2.820 0.560 2.980 1.040 ;
        RECT  0.600 0.560 2.980 0.720 ;
        RECT  2.460 0.880 2.620 2.320 ;
        RECT  2.460 1.380 2.780 1.660 ;
        RECT  2.400 0.880 2.620 1.160 ;
        RECT  1.240 2.150 2.240 2.310 ;
        RECT  2.080 0.920 2.240 2.310 ;
        RECT  2.080 1.460 2.300 1.740 ;
        RECT  1.240 0.920 2.240 1.080 ;
    END
END DFFKHD

MACRO DFFRBCHD
    CLASS CORE ;
    FOREIGN DFFRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.280 1.500 1.850 ;
        RECT  1.180 1.440 1.500 1.720 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.840 9.500 2.390 ;
        RECT  9.280 2.110 9.500 2.390 ;
        RECT  9.280 0.840 9.500 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.240 1.100 8.700 1.300 ;
        RECT  8.500 1.100 8.700 2.090 ;
        RECT  8.240 1.810 8.700 2.090 ;
        RECT  8.240 0.860 8.460 1.300 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.240 -0.280 1.520 0.400 ;
        RECT  6.340 -0.280 6.620 0.400 ;
        RECT  7.280 -0.280 7.560 0.400 ;
        RECT  8.700 -0.280 8.980 0.840 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.800 1.660 3.480 ;
        RECT  5.820 2.800 6.100 3.480 ;
        RECT  6.270 2.800 6.550 3.480 ;
        RECT  5.820 2.860 6.550 3.480 ;
        RECT  8.200 2.800 8.480 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.800 2.600 3.880 2.760 ;
        RECT  3.720 2.140 3.880 2.760 ;
        RECT  5.600 2.480 8.050 2.640 ;
        RECT  7.890 0.440 8.050 2.640 ;
        RECT  2.800 0.460 2.960 2.760 ;
        RECT  5.600 2.140 5.760 2.640 ;
        RECT  7.890 2.300 9.100 2.460 ;
        RECT  8.940 1.300 9.100 2.460 ;
        RECT  2.380 2.300 2.960 2.460 ;
        RECT  3.720 2.140 5.760 2.300 ;
        RECT  2.640 0.460 2.960 0.680 ;
        RECT  7.840 0.440 8.120 0.660 ;
        RECT  6.790 2.160 7.550 2.320 ;
        RECT  7.390 0.980 7.550 2.320 ;
        RECT  7.390 1.460 7.710 1.740 ;
        RECT  3.120 2.220 3.450 2.440 ;
        RECT  3.120 0.440 3.280 2.440 ;
        RECT  7.070 0.620 7.230 1.720 ;
        RECT  6.020 0.620 7.230 0.780 ;
        RECT  6.020 0.440 6.180 0.780 ;
        RECT  3.120 0.440 6.180 0.600 ;
        RECT  5.920 1.820 6.080 2.220 ;
        RECT  4.020 1.820 6.080 1.980 ;
        RECT  5.220 1.080 5.380 1.980 ;
        RECT  5.220 1.080 5.540 1.300 ;
        RECT  3.960 1.080 5.540 1.240 ;
        RECT  3.960 0.840 4.120 1.240 ;
        RECT  5.540 1.460 5.860 1.620 ;
        RECT  5.700 0.760 5.860 1.620 ;
        RECT  4.380 0.760 5.860 0.920 ;
        RECT  5.220 2.460 5.440 2.740 ;
        RECT  4.300 2.460 5.440 2.620 ;
        RECT  3.440 1.400 3.820 1.980 ;
        RECT  3.440 1.400 4.910 1.560 ;
        RECT  3.440 0.840 3.600 1.980 ;
        RECT  0.600 1.710 0.760 2.180 ;
        RECT  2.480 0.880 2.640 2.080 ;
        RECT  0.580 0.440 0.740 1.870 ;
        RECT  2.320 0.520 2.480 1.040 ;
        RECT  0.580 0.560 1.840 0.720 ;
        RECT  1.680 0.520 2.480 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.000 0.840 2.160 2.490 ;
        RECT  2.000 1.380 2.320 1.660 ;
        RECT  0.900 2.380 1.840 2.540 ;
        RECT  1.680 0.920 1.840 2.540 ;
        RECT  0.900 0.920 1.840 1.080 ;
    END
END DFFRBCHD

MACRO DFFRBEHD
    CLASS CORE ;
    FOREIGN DFFRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.280 1.500 1.850 ;
        RECT  1.180 1.440 1.500 1.720 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.840 9.500 2.390 ;
        RECT  9.280 2.110 9.500 2.390 ;
        RECT  9.280 0.840 9.500 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.240 1.840 8.460 2.120 ;
        RECT  8.240 1.040 8.700 1.240 ;
        RECT  8.500 1.040 8.700 2.040 ;
        RECT  8.240 1.840 8.700 2.040 ;
        RECT  8.240 0.960 8.460 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.240 -0.280 1.520 0.400 ;
        RECT  6.340 -0.280 6.620 0.400 ;
        RECT  7.280 -0.280 7.560 0.400 ;
        RECT  8.700 -0.280 8.980 0.580 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.800 1.660 3.480 ;
        RECT  5.820 2.800 6.100 3.480 ;
        RECT  6.270 2.800 6.550 3.480 ;
        RECT  5.820 2.860 6.550 3.480 ;
        RECT  8.700 2.620 8.980 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.800 2.600 3.880 2.760 ;
        RECT  3.720 2.140 3.880 2.760 ;
        RECT  5.600 2.480 8.050 2.640 ;
        RECT  7.890 0.440 8.050 2.640 ;
        RECT  2.800 0.460 2.960 2.760 ;
        RECT  5.600 2.140 5.760 2.640 ;
        RECT  7.890 2.300 9.080 2.460 ;
        RECT  8.920 1.300 9.080 2.460 ;
        RECT  2.380 2.300 2.960 2.460 ;
        RECT  3.720 2.140 5.760 2.300 ;
        RECT  2.640 0.460 2.960 0.680 ;
        RECT  7.840 0.440 8.120 0.660 ;
        RECT  6.790 2.160 7.550 2.320 ;
        RECT  7.390 0.980 7.550 2.320 ;
        RECT  7.390 1.460 7.710 1.740 ;
        RECT  3.120 2.220 3.450 2.440 ;
        RECT  3.120 0.440 3.280 2.440 ;
        RECT  7.070 0.620 7.230 1.720 ;
        RECT  6.020 0.620 7.230 0.780 ;
        RECT  6.020 0.440 6.180 0.780 ;
        RECT  3.120 0.440 6.180 0.600 ;
        RECT  5.920 1.820 6.080 2.220 ;
        RECT  4.020 1.820 6.080 1.980 ;
        RECT  5.220 1.080 5.380 1.980 ;
        RECT  5.220 1.080 5.540 1.300 ;
        RECT  3.960 1.080 5.540 1.240 ;
        RECT  3.960 0.840 4.120 1.240 ;
        RECT  5.540 1.460 5.860 1.620 ;
        RECT  5.700 0.760 5.860 1.620 ;
        RECT  4.380 0.760 5.860 0.920 ;
        RECT  5.220 2.460 5.440 2.740 ;
        RECT  4.300 2.460 5.440 2.620 ;
        RECT  3.440 1.400 3.820 1.980 ;
        RECT  3.440 1.400 4.910 1.560 ;
        RECT  3.440 0.840 3.600 1.980 ;
        RECT  0.600 1.710 0.760 2.180 ;
        RECT  2.480 0.880 2.640 2.080 ;
        RECT  0.580 0.440 0.740 1.870 ;
        RECT  2.320 0.520 2.480 1.040 ;
        RECT  0.580 0.560 1.840 0.720 ;
        RECT  1.680 0.520 2.480 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.000 0.840 2.160 2.340 ;
        RECT  2.000 1.380 2.320 1.660 ;
        RECT  0.900 2.380 1.840 2.540 ;
        RECT  1.680 0.920 1.840 2.540 ;
        RECT  0.900 0.920 1.840 1.080 ;
    END
END DFFRBEHD

MACRO DFFRBHHD
    CLASS CORE ;
    FOREIGN DFFRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.440 1.560 1.720 ;
        RECT  1.300 1.200 1.500 1.740 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.790 10.700 2.360 ;
        RECT  10.360 2.080 10.700 2.360 ;
        RECT  10.360 0.820 10.700 1.100 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.610 9.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.280 1.880 0.400 ;
        RECT  6.610 -0.280 6.890 0.400 ;
        RECT  8.740 -0.280 9.020 0.580 ;
        RECT  9.780 -0.280 10.060 0.580 ;
        RECT  10.820 -0.280 11.100 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.580 2.800 1.860 3.480 ;
        RECT  6.670 2.740 7.010 3.480 ;
        RECT  7.690 2.620 7.970 3.480 ;
        RECT  8.740 2.620 9.020 3.480 ;
        RECT  9.780 2.620 10.060 3.480 ;
        RECT  10.820 2.620 11.100 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.020 2.600 6.510 2.760 ;
        RECT  6.350 2.420 6.510 2.760 ;
        RECT  3.020 0.460 3.180 2.760 ;
        RECT  6.350 2.420 7.480 2.580 ;
        RECT  10.040 1.420 10.200 2.460 ;
        RECT  2.600 2.300 3.180 2.460 ;
        RECT  7.320 2.300 10.200 2.460 ;
        RECT  8.240 0.890 8.400 2.460 ;
        RECT  2.860 0.460 3.180 0.680 ;
        RECT  7.130 1.980 7.850 2.140 ;
        RECT  7.690 0.600 7.850 2.140 ;
        RECT  7.690 1.460 8.050 1.740 ;
        RECT  3.340 2.220 3.670 2.440 ;
        RECT  3.340 0.440 3.500 2.440 ;
        RECT  7.370 0.560 7.530 1.680 ;
        RECT  6.220 0.560 7.530 0.720 ;
        RECT  3.340 0.440 6.380 0.600 ;
        RECT  4.610 2.280 6.190 2.440 ;
        RECT  6.030 1.460 6.190 2.440 ;
        RECT  5.640 1.460 6.190 1.620 ;
        RECT  5.900 0.760 6.060 1.620 ;
        RECT  4.560 0.760 6.060 0.920 ;
        RECT  4.920 1.960 5.870 2.120 ;
        RECT  5.590 1.900 5.870 2.120 ;
        RECT  4.240 1.820 5.080 1.980 ;
        RECT  4.920 1.080 5.080 2.120 ;
        RECT  5.460 1.080 5.740 1.300 ;
        RECT  4.180 1.080 5.740 1.240 ;
        RECT  4.180 0.840 4.340 1.240 ;
        RECT  3.660 1.400 4.040 1.980 ;
        RECT  3.660 1.400 4.750 1.560 ;
        RECT  3.660 0.840 3.820 1.980 ;
        RECT  0.600 1.680 0.760 2.170 ;
        RECT  2.700 0.880 2.860 2.040 ;
        RECT  0.580 0.440 0.740 1.840 ;
        RECT  2.540 0.560 2.700 1.040 ;
        RECT  0.580 0.560 2.700 0.720 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.220 0.880 2.380 2.540 ;
        RECT  2.220 1.380 2.540 1.660 ;
        RECT  2.160 0.880 2.380 1.160 ;
        RECT  0.960 2.420 2.000 2.580 ;
        RECT  1.840 0.880 2.000 2.580 ;
        RECT  1.840 1.440 2.060 1.720 ;
        RECT  0.960 0.880 2.000 1.040 ;
    END
END DFFRBHHD

MACRO DFFRBKHD
    CLASS CORE ;
    FOREIGN DFFRBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.440 1.570 1.720 ;
        RECT  1.300 1.200 1.500 1.740 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.080 0.860 12.770 1.140 ;
        RECT  11.260 2.060 12.770 2.340 ;
        RECT  11.700 0.860 11.900 2.340 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.980 0.860 10.670 1.140 ;
        RECT  8.980 1.840 10.670 2.120 ;
        RECT  9.700 0.860 9.900 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.570 -0.280 1.850 0.400 ;
        RECT  6.620 -0.280 6.900 0.400 ;
        RECT  8.640 -0.280 8.920 0.580 ;
        RECT  9.700 -0.280 9.980 0.580 ;
        RECT  10.740 -0.280 11.020 0.580 ;
        RECT  11.780 -0.280 12.060 0.580 ;
        RECT  12.820 -0.280 13.100 0.580 ;
        RECT  0.000 -0.280 13.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.590 2.800 1.870 3.480 ;
        RECT  6.680 2.740 8.020 3.480 ;
        RECT  8.640 2.620 8.920 3.480 ;
        RECT  9.700 2.620 9.980 3.480 ;
        RECT  10.740 2.620 11.020 3.480 ;
        RECT  11.780 2.620 12.060 3.480 ;
        RECT  12.820 2.620 13.100 3.480 ;
        RECT  0.000 2.920 13.200 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.030 2.600 6.520 2.760 ;
        RECT  6.360 2.420 6.520 2.760 ;
        RECT  3.030 0.460 3.190 2.760 ;
        RECT  6.360 2.420 8.380 2.580 ;
        RECT  8.220 0.890 8.380 2.580 ;
        RECT  10.920 1.460 11.080 2.460 ;
        RECT  2.610 2.300 3.190 2.460 ;
        RECT  8.140 2.300 11.080 2.460 ;
        RECT  8.140 1.840 8.380 2.580 ;
        RECT  10.920 1.460 11.140 1.740 ;
        RECT  8.140 0.890 8.380 1.240 ;
        RECT  2.870 0.460 3.190 0.680 ;
        RECT  7.140 2.100 7.860 2.260 ;
        RECT  7.700 0.770 7.860 2.260 ;
        RECT  7.700 1.400 8.060 1.680 ;
        RECT  7.640 0.770 7.860 1.050 ;
        RECT  3.350 2.220 3.680 2.440 ;
        RECT  3.350 0.440 3.510 2.440 ;
        RECT  7.320 1.400 7.540 1.680 ;
        RECT  7.320 0.560 7.480 1.680 ;
        RECT  6.230 0.560 7.480 0.720 ;
        RECT  3.350 0.440 6.390 0.600 ;
        RECT  4.620 2.280 6.200 2.440 ;
        RECT  6.040 1.460 6.200 2.440 ;
        RECT  5.640 1.460 6.200 1.620 ;
        RECT  5.910 0.760 6.070 1.620 ;
        RECT  4.570 0.760 6.070 0.920 ;
        RECT  4.930 1.960 5.880 2.120 ;
        RECT  5.600 1.900 5.880 2.120 ;
        RECT  4.250 1.820 5.090 1.980 ;
        RECT  4.930 1.080 5.090 2.120 ;
        RECT  5.470 1.080 5.750 1.300 ;
        RECT  4.190 1.080 5.750 1.240 ;
        RECT  4.190 0.840 4.350 1.240 ;
        RECT  3.670 1.400 4.050 1.980 ;
        RECT  3.670 1.400 4.750 1.560 ;
        RECT  3.670 0.840 3.830 1.980 ;
        RECT  0.600 0.440 0.760 2.160 ;
        RECT  2.710 0.880 2.870 2.080 ;
        RECT  2.550 0.520 2.710 1.040 ;
        RECT  0.580 0.560 2.120 0.720 ;
        RECT  1.960 0.520 2.710 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.230 0.840 2.390 2.540 ;
        RECT  2.230 1.380 2.550 1.660 ;
        RECT  0.970 2.360 2.070 2.520 ;
        RECT  1.910 0.880 2.070 2.520 ;
        RECT  0.970 0.880 2.070 1.040 ;
    END
END DFFRBKHD

MACRO DFFRSBEHD
    CLASS CORE ;
    FOREIGN DFFRSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.090 0.840 7.500 1.340 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.420 1.500 1.700 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.480 1.840 10.700 2.120 ;
        RECT  10.500 0.920 10.700 2.160 ;
        RECT  10.480 0.960 10.700 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.320 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 1.020 9.580 1.240 ;
        RECT  9.300 0.980 9.500 2.160 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.420 8.300 1.960 ;
        RECT  8.070 1.420 8.300 1.700 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.310 -0.280 1.590 0.400 ;
        RECT  5.430 -0.280 5.710 0.620 ;
        RECT  6.870 -0.280 7.150 0.620 ;
        RECT  8.090 -0.280 8.370 0.620 ;
        RECT  9.860 -0.280 10.140 0.400 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.470 2.800 1.750 3.480 ;
        RECT  4.930 2.800 5.210 3.480 ;
        RECT  6.530 2.800 6.810 3.480 ;
        RECT  7.690 2.800 7.970 3.480 ;
        RECT  8.710 2.800 8.990 3.480 ;
        RECT  9.860 2.800 10.140 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.890 2.600 4.120 2.760 ;
        RECT  3.960 2.160 4.120 2.760 ;
        RECT  8.820 2.480 10.200 2.640 ;
        RECT  10.040 0.560 10.200 2.640 ;
        RECT  2.890 0.460 3.050 2.760 ;
        RECT  8.820 2.160 8.980 2.640 ;
        RECT  2.510 2.300 3.050 2.460 ;
        RECT  3.960 2.160 8.980 2.320 ;
        RECT  10.040 1.340 10.280 1.620 ;
        RECT  8.930 0.440 9.210 0.750 ;
        RECT  8.930 0.560 10.200 0.720 ;
        RECT  2.730 0.460 3.050 0.680 ;
        RECT  8.870 1.090 9.030 1.750 ;
        RECT  8.440 1.090 9.030 1.250 ;
        RECT  7.750 0.940 8.600 1.100 ;
        RECT  8.220 2.480 8.550 2.740 ;
        RECT  7.050 2.480 8.550 2.640 ;
        RECT  3.520 2.280 3.800 2.440 ;
        RECT  3.560 1.840 3.720 2.440 ;
        RECT  3.560 1.840 4.450 2.000 ;
        RECT  4.290 1.060 4.450 2.000 ;
        RECT  7.490 1.500 7.650 1.920 ;
        RECT  4.290 1.500 7.650 1.660 ;
        RECT  3.870 1.060 4.450 1.220 ;
        RECT  3.870 0.600 4.030 1.220 ;
        RECT  3.250 0.600 4.030 0.760 ;
        RECT  3.250 0.460 3.590 0.760 ;
        RECT  4.610 1.820 7.330 1.980 ;
        RECT  4.280 2.480 6.470 2.640 ;
        RECT  4.720 1.180 6.210 1.340 ;
        RECT  6.050 0.700 6.210 1.340 ;
        RECT  4.720 0.880 4.880 1.340 ;
        RECT  4.610 0.880 4.880 1.160 ;
        RECT  5.040 0.840 5.890 1.000 ;
        RECT  5.040 0.460 5.200 1.000 ;
        RECT  4.220 0.460 5.200 0.620 ;
        RECT  3.210 0.940 3.370 2.080 ;
        RECT  3.210 1.380 4.130 1.660 ;
        RECT  3.210 0.940 3.570 1.100 ;
        RECT  0.610 0.560 0.770 2.230 ;
        RECT  2.570 0.880 2.730 2.040 ;
        RECT  2.410 0.440 2.570 1.040 ;
        RECT  0.610 0.560 1.910 0.720 ;
        RECT  1.750 0.440 2.570 0.600 ;
        RECT  2.090 0.760 2.250 2.340 ;
        RECT  2.090 1.380 2.390 1.660 ;
        RECT  1.030 2.180 1.910 2.340 ;
        RECT  1.750 0.880 1.910 2.340 ;
        RECT  1.030 0.880 1.910 1.040 ;
    END
END DFFRSBEHD

MACRO DFFRSBHHD
    CLASS CORE ;
    FOREIGN DFFRSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 1.640 7.500 2.140 ;
        RECT  7.280 1.780 7.500 2.060 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.420 1.500 1.700 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.920 11.500 2.160 ;
        RECT  11.160 1.840 11.500 2.160 ;
        RECT  11.160 0.920 11.500 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.320 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.060 0.960 10.340 1.240 ;
        RECT  10.060 1.840 10.340 2.120 ;
        RECT  10.100 0.960 10.300 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.420 8.700 1.960 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.310 -0.280 1.590 0.400 ;
        RECT  5.480 -0.280 5.700 0.680 ;
        RECT  7.000 -0.280 7.280 0.620 ;
        RECT  8.320 -0.280 8.600 0.620 ;
        RECT  9.500 -0.280 9.780 0.400 ;
        RECT  10.580 -0.280 10.860 0.580 ;
        RECT  11.620 -0.280 11.900 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.470 2.800 1.750 3.480 ;
        RECT  4.930 2.800 5.210 3.480 ;
        RECT  6.350 2.800 6.630 3.480 ;
        RECT  7.180 2.800 7.460 3.480 ;
        RECT  8.380 2.800 8.660 3.480 ;
        RECT  9.500 2.800 9.780 3.480 ;
        RECT  10.580 2.620 10.860 3.480 ;
        RECT  11.620 2.620 11.900 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.890 2.600 4.120 2.760 ;
        RECT  3.960 2.160 4.120 2.760 ;
        RECT  6.450 2.480 10.350 2.640 ;
        RECT  10.190 2.280 10.350 2.640 ;
        RECT  2.890 0.460 3.050 2.760 ;
        RECT  9.720 0.900 9.880 2.640 ;
        RECT  6.450 2.160 6.610 2.640 ;
        RECT  2.510 2.300 3.050 2.460 ;
        RECT  10.190 2.280 11.000 2.440 ;
        RECT  10.840 1.300 11.000 2.440 ;
        RECT  3.960 2.160 6.610 2.320 ;
        RECT  9.220 0.900 9.880 1.060 ;
        RECT  9.220 0.750 9.440 1.060 ;
        RECT  2.730 0.460 3.050 0.680 ;
        RECT  7.740 2.160 9.480 2.320 ;
        RECT  9.320 1.240 9.480 2.320 ;
        RECT  8.880 1.240 9.480 1.400 ;
        RECT  8.880 0.780 9.040 1.400 ;
        RECT  7.840 0.780 8.160 1.040 ;
        RECT  7.840 0.780 9.040 0.940 ;
        RECT  3.520 2.280 3.800 2.440 ;
        RECT  3.560 1.840 3.720 2.440 ;
        RECT  3.560 1.840 4.450 2.000 ;
        RECT  4.290 1.060 4.450 2.000 ;
        RECT  8.060 1.200 8.220 1.940 ;
        RECT  4.290 1.500 6.770 1.660 ;
        RECT  6.610 1.200 6.770 1.660 ;
        RECT  6.610 1.200 8.220 1.360 ;
        RECT  3.870 1.060 4.450 1.220 ;
        RECT  3.870 0.600 4.030 1.220 ;
        RECT  3.250 0.600 4.030 0.760 ;
        RECT  3.250 0.460 3.590 0.760 ;
        RECT  6.770 2.100 7.110 2.320 ;
        RECT  6.770 1.820 6.930 2.320 ;
        RECT  4.610 1.820 6.930 1.980 ;
        RECT  5.040 0.840 6.020 1.000 ;
        RECT  5.860 0.560 6.020 1.000 ;
        RECT  5.040 0.460 5.200 1.000 ;
        RECT  5.860 0.560 6.580 0.720 ;
        RECT  4.220 0.460 5.200 0.620 ;
        RECT  4.720 1.180 6.400 1.340 ;
        RECT  6.180 0.880 6.400 1.340 ;
        RECT  4.720 0.880 4.880 1.340 ;
        RECT  4.610 0.880 4.880 1.160 ;
        RECT  4.280 2.480 6.290 2.640 ;
        RECT  3.210 0.940 3.370 2.080 ;
        RECT  3.210 1.380 4.130 1.660 ;
        RECT  3.210 0.940 3.570 1.100 ;
        RECT  0.610 0.560 0.770 2.230 ;
        RECT  2.570 0.880 2.730 2.040 ;
        RECT  2.410 0.440 2.570 1.040 ;
        RECT  0.610 0.560 1.910 0.720 ;
        RECT  1.750 0.440 2.570 0.600 ;
        RECT  2.090 0.760 2.250 2.340 ;
        RECT  2.090 1.380 2.390 1.660 ;
        RECT  1.030 2.180 1.910 2.340 ;
        RECT  1.750 0.880 1.910 2.340 ;
        RECT  1.030 0.880 1.910 1.040 ;
    END
END DFFRSBHHD

MACRO DFFSBEHD
    CLASS CORE ;
    FOREIGN DFFSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.480 1.500 1.760 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.840 9.500 2.260 ;
        RECT  9.270 1.980 9.500 2.260 ;
        RECT  9.270 0.840 9.500 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.980 8.700 2.140 ;
        RECT  8.170 1.940 8.700 2.140 ;
        RECT  8.170 0.980 8.700 1.180 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.140 6.300 1.660 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.580 0.400 ;
        RECT  4.980 -0.280 5.260 0.400 ;
        RECT  7.690 -0.280 7.970 0.400 ;
        RECT  8.690 -0.280 8.970 0.580 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 2.800 1.740 3.480 ;
        RECT  4.970 2.800 5.250 3.480 ;
        RECT  5.730 2.800 6.010 3.480 ;
        RECT  6.970 2.800 7.250 3.480 ;
        RECT  8.690 2.620 8.970 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.880 2.600 3.870 2.760 ;
        RECT  3.710 2.160 3.870 2.760 ;
        RECT  4.850 2.480 8.390 2.640 ;
        RECT  8.230 2.300 8.390 2.640 ;
        RECT  2.880 0.460 3.040 2.760 ;
        RECT  6.730 0.940 6.890 2.640 ;
        RECT  4.850 2.160 5.010 2.640 ;
        RECT  8.230 2.300 9.090 2.460 ;
        RECT  8.930 1.460 9.090 2.460 ;
        RECT  2.500 2.300 3.040 2.460 ;
        RECT  3.710 2.160 5.010 2.320 ;
        RECT  8.930 1.460 9.140 1.740 ;
        RECT  6.730 0.940 7.210 1.100 ;
        RECT  2.720 0.460 3.040 0.680 ;
        RECT  7.690 2.100 7.970 2.260 ;
        RECT  7.690 1.780 7.910 2.260 ;
        RECT  7.750 0.700 7.910 2.260 ;
        RECT  7.090 1.780 7.910 1.940 ;
        RECT  7.090 1.620 7.250 1.940 ;
        RECT  7.750 1.410 8.340 1.690 ;
        RECT  3.200 2.280 3.550 2.440 ;
        RECT  3.200 0.460 3.360 2.440 ;
        RECT  7.370 0.440 7.530 1.400 ;
        RECT  3.840 0.990 5.080 1.150 ;
        RECT  4.920 0.560 5.080 1.150 ;
        RECT  3.840 0.460 4.000 1.150 ;
        RECT  4.920 0.560 5.620 0.720 ;
        RECT  3.200 0.460 4.000 0.620 ;
        RECT  5.460 0.440 7.530 0.600 ;
        RECT  5.250 2.160 5.720 2.320 ;
        RECT  5.560 1.340 5.720 2.320 ;
        RECT  5.560 1.920 6.570 2.080 ;
        RECT  4.310 1.340 5.720 1.500 ;
        RECT  5.290 0.940 5.570 1.500 ;
        RECT  3.520 1.820 5.400 1.980 ;
        RECT  5.120 1.680 5.400 1.980 ;
        RECT  3.520 0.840 3.680 1.980 ;
        RECT  4.160 0.460 4.760 0.740 ;
        RECT  4.030 2.480 4.570 2.760 ;
        RECT  0.600 0.560 0.760 2.230 ;
        RECT  2.560 0.880 2.720 2.040 ;
        RECT  2.400 0.440 2.560 1.040 ;
        RECT  0.600 0.560 1.900 0.720 ;
        RECT  1.740 0.440 2.560 0.600 ;
        RECT  2.080 0.760 2.240 2.400 ;
        RECT  2.080 1.380 2.380 1.660 ;
        RECT  1.020 2.180 1.900 2.340 ;
        RECT  1.740 0.910 1.900 2.340 ;
        RECT  1.020 0.910 1.900 1.070 ;
    END
END DFFSBEHD

MACRO DFFSBHHD
    CLASS CORE ;
    FOREIGN DFFSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.480 1.500 1.760 ;
        END
    END CK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.800 10.700 2.360 ;
        RECT  10.360 2.080 10.700 2.360 ;
        RECT  10.360 0.800 10.700 1.080 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.800 9.500 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.380 6.350 1.660 ;
        RECT  6.100 1.140 6.300 1.660 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.580 0.400 ;
        RECT  4.990 -0.280 5.270 0.400 ;
        RECT  6.470 -0.280 6.750 0.400 ;
        RECT  8.700 -0.280 8.980 0.400 ;
        RECT  9.780 -0.280 10.060 0.580 ;
        RECT  10.820 -0.280 11.100 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 2.800 1.740 3.480 ;
        RECT  5.010 2.800 6.140 3.480 ;
        RECT  6.700 2.800 6.980 3.480 ;
        RECT  7.820 2.800 8.100 3.480 ;
        RECT  8.740 2.620 9.020 3.480 ;
        RECT  9.780 2.620 10.060 3.480 ;
        RECT  10.820 2.620 11.100 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.880 2.600 3.870 2.760 ;
        RECT  3.710 2.160 3.870 2.760 ;
        RECT  4.950 2.480 7.480 2.640 ;
        RECT  7.320 1.020 7.480 2.640 ;
        RECT  2.880 0.460 3.040 2.760 ;
        RECT  4.950 2.160 5.110 2.640 ;
        RECT  2.500 2.300 3.040 2.460 ;
        RECT  7.320 2.280 10.200 2.440 ;
        RECT  10.040 1.400 10.200 2.440 ;
        RECT  3.710 2.160 5.110 2.320 ;
        RECT  7.320 1.020 7.740 1.180 ;
        RECT  2.720 0.460 3.040 0.680 ;
        RECT  8.180 1.960 9.140 2.120 ;
        RECT  8.980 1.400 9.140 2.120 ;
        RECT  8.180 0.960 8.340 2.120 ;
        RECT  8.020 0.960 8.340 1.620 ;
        RECT  3.200 2.280 3.550 2.440 ;
        RECT  3.200 0.460 3.360 2.440 ;
        RECT  8.500 0.640 8.660 1.620 ;
        RECT  3.840 0.990 5.250 1.150 ;
        RECT  5.090 0.560 5.250 1.150 ;
        RECT  3.840 0.460 4.000 1.150 ;
        RECT  8.200 0.640 8.660 0.800 ;
        RECT  5.090 0.560 8.360 0.720 ;
        RECT  3.200 0.460 4.000 0.620 ;
        RECT  5.270 2.160 5.750 2.320 ;
        RECT  5.590 0.940 5.750 2.320 ;
        RECT  5.590 2.100 6.630 2.260 ;
        RECT  4.410 1.340 5.750 1.500 ;
        RECT  5.470 0.940 5.750 1.500 ;
        RECT  3.520 1.820 5.400 1.980 ;
        RECT  5.080 1.660 5.400 1.980 ;
        RECT  3.520 0.840 3.680 1.980 ;
        RECT  4.250 2.480 4.790 2.760 ;
        RECT  4.160 0.460 4.780 0.740 ;
        RECT  0.600 0.560 0.760 2.230 ;
        RECT  2.560 0.880 2.720 2.040 ;
        RECT  2.400 0.440 2.560 1.040 ;
        RECT  0.600 0.560 1.900 0.720 ;
        RECT  1.740 0.440 2.560 0.600 ;
        RECT  2.080 0.760 2.240 2.400 ;
        RECT  2.080 1.380 2.380 1.660 ;
        RECT  1.020 2.180 1.900 2.340 ;
        RECT  1.740 0.910 1.900 2.340 ;
        RECT  1.020 0.910 1.900 1.070 ;
    END
END DFFSBHHD

MACRO DFTRBCHD
    CLASS CORE ;
    FOREIGN DFTRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.870 9.900 2.160 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.910 ;
        RECT  1.180 1.410 1.500 1.690 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.840 10.700 1.560 ;
        RECT  10.480 1.140 10.700 1.420 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.340 2.100 8.540 2.720 ;
        RECT  8.500 0.960 8.700 2.300 ;
        RECT  8.300 0.960 8.700 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  6.340 -0.280 6.620 0.400 ;
        RECT  7.330 -0.280 7.610 0.400 ;
        RECT  8.800 -0.280 9.080 0.580 ;
        RECT  10.120 -0.280 10.400 0.400 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.800 1.660 3.480 ;
        RECT  5.820 2.800 6.550 3.480 ;
        RECT  7.390 2.800 7.670 3.480 ;
        RECT  8.800 2.620 9.080 3.480 ;
        RECT  10.150 2.800 10.430 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.120 1.620 10.340 2.500 ;
        RECT  10.120 0.700 10.280 2.500 ;
        RECT  10.120 0.700 10.340 0.980 ;
        RECT  2.800 2.600 3.880 2.760 ;
        RECT  3.720 2.140 3.880 2.760 ;
        RECT  5.600 2.480 8.050 2.640 ;
        RECT  7.890 0.460 8.050 2.640 ;
        RECT  2.800 0.460 2.960 2.760 ;
        RECT  5.600 2.140 5.760 2.640 ;
        RECT  2.380 2.300 2.960 2.460 ;
        RECT  3.720 2.140 5.760 2.300 ;
        RECT  7.890 0.460 8.120 0.740 ;
        RECT  2.640 0.460 2.960 0.680 ;
        RECT  6.790 2.160 7.550 2.320 ;
        RECT  7.390 0.980 7.550 2.320 ;
        RECT  7.390 1.460 7.710 1.740 ;
        RECT  3.120 2.220 3.450 2.440 ;
        RECT  3.120 0.440 3.280 2.440 ;
        RECT  7.070 0.620 7.230 1.720 ;
        RECT  6.020 0.620 7.230 0.780 ;
        RECT  6.020 0.440 6.180 0.780 ;
        RECT  3.120 0.440 6.180 0.600 ;
        RECT  5.920 1.820 6.080 2.230 ;
        RECT  4.020 1.820 6.080 1.980 ;
        RECT  5.100 1.080 5.260 1.980 ;
        RECT  5.100 1.080 5.540 1.300 ;
        RECT  3.960 1.080 5.540 1.240 ;
        RECT  3.960 0.840 4.120 1.240 ;
        RECT  5.540 1.460 5.860 1.620 ;
        RECT  5.700 0.760 5.860 1.620 ;
        RECT  4.340 0.760 5.860 0.920 ;
        RECT  5.220 2.460 5.440 2.740 ;
        RECT  4.300 2.460 5.440 2.620 ;
        RECT  3.440 1.400 3.820 1.980 ;
        RECT  3.440 1.400 4.900 1.560 ;
        RECT  3.440 0.840 3.600 1.980 ;
        RECT  0.540 1.840 0.760 2.120 ;
        RECT  2.480 0.880 2.640 2.080 ;
        RECT  0.580 0.440 0.740 2.120 ;
        RECT  2.320 0.520 2.480 1.040 ;
        RECT  0.580 0.560 1.890 0.720 ;
        RECT  1.730 0.520 2.480 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.000 0.840 2.160 2.440 ;
        RECT  2.000 1.380 2.320 1.660 ;
        RECT  0.860 2.370 1.840 2.530 ;
        RECT  1.680 0.910 1.840 2.530 ;
        RECT  0.900 0.910 1.840 1.070 ;
    END
END DFTRBCHD

MACRO DFTRBEHD
    CLASS CORE ;
    FOREIGN DFTRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.840 11.100 2.360 ;
        RECT  10.740 2.060 11.100 2.360 ;
        RECT  10.740 0.840 11.100 1.140 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.910 ;
        RECT  1.180 1.410 1.500 1.690 ;
        END
    END CK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.100 1.140 12.300 1.860 ;
        RECT  12.080 1.140 12.300 1.420 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.960 8.700 2.120 ;
        RECT  8.380 1.840 8.700 2.120 ;
        RECT  8.380 0.960 8.700 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.370 -0.280 1.650 0.400 ;
        RECT  6.370 -0.280 6.650 0.400 ;
        RECT  7.420 -0.280 7.700 0.400 ;
        RECT  8.840 -0.280 9.120 0.580 ;
        RECT  9.880 -0.280 10.160 0.580 ;
        RECT  11.800 -0.280 12.080 0.400 ;
        RECT  0.000 -0.280 12.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 2.800 1.690 3.480 ;
        RECT  5.850 2.800 6.580 3.480 ;
        RECT  7.420 2.800 7.700 3.480 ;
        RECT  8.840 2.620 9.120 3.480 ;
        RECT  9.880 2.620 10.160 3.480 ;
        RECT  11.770 2.800 12.050 3.480 ;
        RECT  0.000 2.920 12.400 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.720 2.000 11.960 2.280 ;
        RECT  11.720 0.800 11.880 2.280 ;
        RECT  11.720 0.800 12.020 0.960 ;
        RECT  11.320 0.520 11.480 1.130 ;
        RECT  9.310 0.920 10.500 1.080 ;
        RECT  10.340 0.520 10.500 1.080 ;
        RECT  10.340 0.520 11.480 0.680 ;
        RECT  10.340 2.520 11.480 2.680 ;
        RECT  11.320 2.050 11.480 2.680 ;
        RECT  10.340 2.120 10.500 2.680 ;
        RECT  9.310 2.120 10.500 2.280 ;
        RECT  2.830 2.600 3.910 2.760 ;
        RECT  3.750 2.140 3.910 2.760 ;
        RECT  5.630 2.480 8.200 2.640 ;
        RECT  8.040 0.480 8.200 2.640 ;
        RECT  2.830 0.460 2.990 2.760 ;
        RECT  5.630 2.140 5.790 2.640 ;
        RECT  2.410 2.300 2.990 2.460 ;
        RECT  3.750 2.140 5.790 2.300 ;
        RECT  7.980 0.480 8.200 0.760 ;
        RECT  2.670 0.460 2.990 0.680 ;
        RECT  6.820 2.160 7.580 2.320 ;
        RECT  7.420 0.980 7.580 2.320 ;
        RECT  7.420 1.460 7.740 1.740 ;
        RECT  3.150 2.220 3.480 2.440 ;
        RECT  3.150 0.440 3.310 2.440 ;
        RECT  7.100 0.620 7.260 1.720 ;
        RECT  6.050 0.620 7.260 0.780 ;
        RECT  6.050 0.440 6.210 0.780 ;
        RECT  3.150 0.440 6.210 0.600 ;
        RECT  5.950 1.820 6.110 2.230 ;
        RECT  4.050 1.820 6.110 1.980 ;
        RECT  5.130 1.080 5.290 1.980 ;
        RECT  5.130 1.080 5.570 1.300 ;
        RECT  3.990 1.080 5.570 1.240 ;
        RECT  3.990 0.840 4.150 1.240 ;
        RECT  5.570 1.460 5.890 1.620 ;
        RECT  5.730 0.760 5.890 1.620 ;
        RECT  4.370 0.760 5.890 0.920 ;
        RECT  5.250 2.460 5.470 2.740 ;
        RECT  4.330 2.460 5.470 2.620 ;
        RECT  3.470 1.400 3.850 1.980 ;
        RECT  3.470 1.400 4.930 1.560 ;
        RECT  3.470 0.840 3.630 1.980 ;
        RECT  0.540 1.840 0.760 2.120 ;
        RECT  2.510 0.880 2.670 2.080 ;
        RECT  0.580 0.440 0.740 2.120 ;
        RECT  2.350 0.520 2.510 1.040 ;
        RECT  0.580 0.560 1.920 0.720 ;
        RECT  1.760 0.520 2.510 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.030 0.840 2.190 2.440 ;
        RECT  2.030 1.380 2.350 1.660 ;
        RECT  0.890 2.350 1.870 2.510 ;
        RECT  1.710 0.900 1.870 2.510 ;
        RECT  0.930 0.900 1.870 1.060 ;
    END
END DFTRBEHD

MACRO DFZCHD
    CLASS CORE ;
    FOREIGN DFZCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.310 3.190 1.590 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 0.580 10.300 2.120 ;
        RECT  10.080 1.840 10.300 2.120 ;
        RECT  10.080 0.580 10.300 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.300 9.100 2.120 ;
        RECT  9.060 0.440 9.260 1.500 ;
        RECT  8.880 0.440 9.260 0.600 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 3.420 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  8.180 -0.280 8.460 0.420 ;
        RECT  9.560 -0.280 9.780 0.660 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.520 3.480 ;
        RECT  6.570 2.800 6.850 3.480 ;
        RECT  7.620 2.800 8.360 3.480 ;
        RECT  9.540 2.800 9.820 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  8.580 2.480 8.920 2.720 ;
        RECT  7.710 2.480 9.880 2.640 ;
        RECT  9.720 1.210 9.880 2.640 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  8.580 0.860 8.740 2.720 ;
        RECT  7.710 1.860 7.870 2.640 ;
        RECT  4.240 2.300 4.820 2.460 ;
        RECT  5.490 2.160 6.030 2.320 ;
        RECT  5.870 1.860 6.030 2.320 ;
        RECT  5.870 1.860 7.870 2.020 ;
        RECT  8.570 0.860 8.900 1.080 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  8.120 0.580 8.280 2.120 ;
        RECT  8.120 1.340 8.420 1.620 ;
        RECT  7.580 0.580 8.280 0.740 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.780 1.140 7.940 1.660 ;
        RECT  5.620 1.140 7.940 1.300 ;
        RECT  5.620 0.460 5.780 1.300 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  7.140 0.580 7.420 0.980 ;
        RECT  5.940 0.580 7.420 0.740 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  5.900 2.480 6.430 2.640 ;
        RECT  7.140 2.180 7.420 2.520 ;
        RECT  6.270 2.360 7.420 2.520 ;
        RECT  5.300 1.460 5.700 1.980 ;
        RECT  5.300 1.460 7.280 1.620 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.660 0.560 3.740 0.720 ;
        RECT  3.580 0.440 4.380 0.600 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  3.860 0.840 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.920 3.680 2.310 ;
        RECT  2.760 0.920 3.680 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END DFZCHD

MACRO DFZCLRBEHD
    CLASS CORE ;
    FOREIGN DFZCLRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.120 1.740 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.350 8.390 1.630 ;
        RECT  8.100 1.240 8.300 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 1.460 7.200 1.740 ;
        RECT  6.900 1.140 7.100 1.790 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.300 0.580 15.500 2.120 ;
        RECT  15.280 1.840 15.500 2.120 ;
        RECT  15.280 0.580 15.500 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 1.900 2.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.100 1.300 14.300 2.120 ;
        RECT  14.260 0.440 14.460 1.500 ;
        RECT  14.180 0.440 14.460 0.660 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.350 5.240 1.630 ;
        RECT  4.900 1.120 5.100 1.680 ;
        END
    END SEL
    PIN LD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.820 0.700 2.640 ;
        RECT  0.500 2.480 2.980 2.640 ;
        RECT  2.820 2.600 3.940 2.760 ;
        RECT  0.480 1.820 0.700 2.100 ;
        END
    END LD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.360 -0.280 4.640 0.400 ;
        RECT  5.000 -0.280 5.280 0.400 ;
        RECT  6.520 -0.280 6.800 0.620 ;
        RECT  8.250 -0.280 8.530 0.400 ;
        RECT  11.900 -0.280 12.180 0.420 ;
        RECT  13.380 -0.280 13.660 0.420 ;
        RECT  14.760 -0.280 14.980 0.660 ;
        RECT  0.000 -0.280 15.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 2.800 2.660 3.480 ;
        RECT  4.440 2.800 5.400 3.480 ;
        RECT  7.080 2.800 7.360 3.480 ;
        RECT  8.440 2.800 8.720 3.480 ;
        RECT  11.770 2.800 12.050 3.480 ;
        RECT  12.820 2.800 13.560 3.480 ;
        RECT  14.700 2.620 14.980 3.480 ;
        RECT  0.000 2.920 15.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.860 2.600 10.850 2.760 ;
        RECT  10.690 2.160 10.850 2.760 ;
        RECT  13.780 2.300 14.120 2.720 ;
        RECT  12.910 2.480 14.120 2.640 ;
        RECT  9.480 2.300 10.020 2.640 ;
        RECT  4.260 2.480 10.020 2.640 ;
        RECT  12.910 1.860 13.070 2.640 ;
        RECT  4.260 2.280 4.420 2.640 ;
        RECT  13.780 2.300 15.080 2.460 ;
        RECT  14.920 1.210 15.080 2.460 ;
        RECT  3.140 2.280 4.420 2.440 ;
        RECT  10.690 2.160 11.230 2.320 ;
        RECT  11.070 1.860 11.230 2.320 ;
        RECT  13.780 0.860 13.940 2.720 ;
        RECT  9.860 0.460 10.020 2.760 ;
        RECT  3.140 1.240 3.300 2.440 ;
        RECT  11.070 1.860 13.070 2.020 ;
        RECT  2.870 1.240 3.300 1.460 ;
        RECT  13.770 0.860 14.100 1.080 ;
        RECT  9.740 0.460 10.020 0.680 ;
        RECT  13.320 0.580 13.480 2.080 ;
        RECT  13.320 1.340 13.620 1.620 ;
        RECT  12.780 0.580 13.480 0.740 ;
        RECT  10.180 2.180 10.530 2.440 ;
        RECT  10.180 0.460 10.340 2.440 ;
        RECT  12.980 1.140 13.140 1.660 ;
        RECT  10.820 1.140 13.140 1.300 ;
        RECT  10.820 0.460 10.980 1.300 ;
        RECT  10.180 0.460 10.980 0.620 ;
        RECT  12.340 0.580 12.620 0.980 ;
        RECT  11.140 0.580 12.620 0.740 ;
        RECT  11.140 0.460 11.740 0.740 ;
        RECT  11.100 2.480 11.630 2.640 ;
        RECT  12.340 2.180 12.620 2.520 ;
        RECT  11.470 2.360 12.620 2.520 ;
        RECT  10.500 1.460 10.900 1.980 ;
        RECT  10.500 1.460 12.480 1.620 ;
        RECT  10.500 0.840 10.660 1.980 ;
        RECT  6.160 2.160 7.620 2.320 ;
        RECT  7.460 0.560 7.620 2.320 ;
        RECT  9.540 0.880 9.700 2.080 ;
        RECT  9.420 0.440 9.580 1.040 ;
        RECT  6.200 0.780 7.620 0.940 ;
        RECT  6.200 0.460 6.360 0.940 ;
        RECT  7.460 0.560 8.880 0.720 ;
        RECT  5.560 0.460 6.360 0.620 ;
        RECT  8.720 0.440 9.580 0.600 ;
        RECT  9.060 0.760 9.220 2.320 ;
        RECT  9.060 1.380 9.360 1.660 ;
        RECT  7.960 2.150 8.880 2.310 ;
        RECT  8.720 0.920 8.880 2.310 ;
        RECT  7.960 0.920 8.880 1.080 ;
        RECT  4.700 2.160 5.980 2.320 ;
        RECT  5.820 1.840 5.980 2.320 ;
        RECT  5.820 1.840 6.560 2.000 ;
        RECT  6.400 1.120 6.560 2.000 ;
        RECT  5.860 1.120 6.560 1.280 ;
        RECT  5.860 0.780 6.020 1.280 ;
        RECT  4.960 0.780 6.020 0.940 ;
        RECT  3.940 1.840 4.480 2.120 ;
        RECT  3.940 1.840 5.660 2.000 ;
        RECT  5.500 1.520 5.660 2.000 ;
        RECT  4.120 0.600 4.280 2.120 ;
        RECT  5.500 1.520 6.140 1.680 ;
        RECT  3.760 0.600 4.280 0.760 ;
        RECT  1.330 2.160 2.710 2.320 ;
        RECT  2.550 0.780 2.710 2.320 ;
        RECT  3.460 1.340 3.680 2.120 ;
        RECT  3.460 1.340 3.920 1.620 ;
        RECT  3.460 0.880 3.620 2.120 ;
        RECT  3.020 0.880 3.620 1.040 ;
        RECT  1.980 0.780 3.180 0.940 ;
        RECT  1.180 0.680 1.460 0.900 ;
        RECT  1.300 0.460 1.460 0.900 ;
        RECT  1.300 0.460 3.180 0.620 ;
        RECT  0.160 0.910 0.320 2.520 ;
        RECT  2.220 1.100 2.380 1.560 ;
        RECT  0.160 1.100 2.380 1.260 ;
    END
END DFZCLRBEHD

MACRO DFZCLRBHHD
    CLASS CORE ;
    FOREIGN DFZCLRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.120 1.740 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.350 8.390 1.630 ;
        RECT  8.100 1.240 8.300 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 1.460 7.200 1.740 ;
        RECT  6.900 1.140 7.100 1.790 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.100 0.840 16.300 2.360 ;
        RECT  15.960 2.080 16.300 2.360 ;
        RECT  15.960 0.840 16.300 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 1.900 2.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.900 0.960 15.100 2.260 ;
        RECT  14.840 1.980 15.100 2.260 ;
        RECT  14.840 0.960 15.100 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.350 5.240 1.630 ;
        RECT  4.900 1.120 5.100 1.680 ;
        END
    END SEL
    PIN LD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.820 0.700 2.640 ;
        RECT  0.500 2.480 2.980 2.640 ;
        RECT  2.820 2.600 3.940 2.760 ;
        RECT  0.480 1.820 0.700 2.100 ;
        END
    END LD
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.360 -0.280 4.640 0.400 ;
        RECT  5.000 -0.280 5.280 0.400 ;
        RECT  6.520 -0.280 6.800 0.620 ;
        RECT  8.250 -0.280 8.530 0.400 ;
        RECT  11.900 -0.280 12.180 0.420 ;
        RECT  12.760 -0.280 13.040 0.420 ;
        RECT  14.220 -0.280 14.500 0.400 ;
        RECT  15.340 -0.280 15.620 0.400 ;
        RECT  16.420 -0.280 16.700 0.580 ;
        RECT  0.000 -0.280 16.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 2.800 2.660 3.480 ;
        RECT  4.440 2.800 5.400 3.480 ;
        RECT  7.080 2.800 7.360 3.480 ;
        RECT  8.440 2.800 8.720 3.480 ;
        RECT  11.770 2.800 12.050 3.480 ;
        RECT  12.760 2.800 13.040 3.480 ;
        RECT  14.220 2.800 14.500 3.480 ;
        RECT  15.340 2.800 15.620 3.480 ;
        RECT  16.420 2.620 16.700 3.480 ;
        RECT  0.000 2.920 16.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.860 2.600 10.850 2.760 ;
        RECT  10.690 2.160 10.850 2.760 ;
        RECT  12.860 2.480 15.800 2.640 ;
        RECT  15.640 0.560 15.800 2.640 ;
        RECT  9.480 2.300 10.020 2.640 ;
        RECT  4.260 2.480 10.020 2.640 ;
        RECT  12.860 1.860 13.020 2.640 ;
        RECT  4.260 2.280 4.420 2.640 ;
        RECT  3.140 2.280 4.420 2.440 ;
        RECT  10.690 2.160 11.230 2.320 ;
        RECT  11.070 1.860 11.230 2.320 ;
        RECT  9.860 0.460 10.020 2.760 ;
        RECT  3.140 1.240 3.300 2.440 ;
        RECT  11.070 1.860 13.020 2.020 ;
        RECT  2.870 1.240 3.300 1.460 ;
        RECT  13.660 0.540 13.940 0.760 ;
        RECT  13.660 0.560 15.800 0.720 ;
        RECT  9.740 0.460 10.020 0.680 ;
        RECT  13.260 1.840 13.540 2.120 ;
        RECT  13.260 0.960 13.420 2.120 ;
        RECT  13.260 1.480 14.320 1.640 ;
        RECT  13.260 0.960 13.540 1.240 ;
        RECT  10.180 2.180 10.530 2.440 ;
        RECT  10.180 0.460 10.340 2.440 ;
        RECT  12.920 1.140 13.080 1.690 ;
        RECT  10.820 1.140 13.080 1.300 ;
        RECT  10.820 0.460 10.980 1.300 ;
        RECT  10.180 0.460 10.980 0.620 ;
        RECT  12.340 0.580 12.620 0.980 ;
        RECT  11.140 0.580 12.620 0.740 ;
        RECT  11.140 0.460 11.740 0.740 ;
        RECT  11.100 2.480 11.630 2.640 ;
        RECT  12.340 2.180 12.620 2.520 ;
        RECT  11.470 2.360 12.620 2.520 ;
        RECT  10.500 1.460 10.900 1.980 ;
        RECT  10.500 1.460 12.480 1.620 ;
        RECT  10.500 0.840 10.660 1.980 ;
        RECT  6.160 2.160 7.620 2.320 ;
        RECT  7.460 0.560 7.620 2.320 ;
        RECT  9.540 0.880 9.700 2.080 ;
        RECT  9.420 0.440 9.580 1.040 ;
        RECT  6.200 0.780 7.620 0.940 ;
        RECT  6.200 0.460 6.360 0.940 ;
        RECT  7.460 0.560 8.880 0.720 ;
        RECT  5.560 0.460 6.360 0.620 ;
        RECT  8.720 0.440 9.580 0.600 ;
        RECT  9.060 0.760 9.220 2.320 ;
        RECT  9.060 1.380 9.360 1.660 ;
        RECT  7.960 2.150 8.880 2.310 ;
        RECT  8.720 0.920 8.880 2.310 ;
        RECT  7.960 0.920 8.880 1.080 ;
        RECT  4.700 2.160 5.980 2.320 ;
        RECT  5.820 1.840 5.980 2.320 ;
        RECT  5.820 1.840 6.560 2.000 ;
        RECT  6.400 1.120 6.560 2.000 ;
        RECT  5.860 1.120 6.560 1.280 ;
        RECT  5.860 0.780 6.020 1.280 ;
        RECT  4.960 0.780 6.020 0.940 ;
        RECT  3.940 1.840 4.480 2.120 ;
        RECT  3.940 1.840 5.660 2.000 ;
        RECT  5.500 1.520 5.660 2.000 ;
        RECT  4.120 0.600 4.280 2.120 ;
        RECT  5.500 1.520 6.140 1.680 ;
        RECT  3.760 0.600 4.280 0.760 ;
        RECT  1.330 2.160 2.710 2.320 ;
        RECT  2.550 0.780 2.710 2.320 ;
        RECT  3.460 1.340 3.680 2.120 ;
        RECT  3.460 1.340 3.920 1.620 ;
        RECT  3.460 0.880 3.620 2.120 ;
        RECT  3.020 0.880 3.620 1.040 ;
        RECT  1.980 0.780 3.180 0.940 ;
        RECT  1.180 0.680 1.460 0.900 ;
        RECT  1.300 0.460 1.460 0.900 ;
        RECT  1.300 0.460 3.180 0.620 ;
        RECT  0.160 0.910 0.320 2.520 ;
        RECT  2.220 1.100 2.380 1.560 ;
        RECT  0.160 1.100 2.380 1.260 ;
    END
END DFZCLRBHHD

MACRO DFZCRBEHD
    CLASS CORE ;
    FOREIGN DFZCRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.420 1.900 2.000 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.350 4.010 1.630 ;
        RECT  3.700 1.240 3.900 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.890 3.500 2.460 ;
        RECT  3.290 1.900 3.500 2.180 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.580 11.100 2.120 ;
        RECT  10.880 1.840 11.100 2.120 ;
        RECT  10.880 0.580 11.100 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 2.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.880 0.440 10.080 1.100 ;
        RECT  9.880 0.900 10.300 1.100 ;
        RECT  10.100 0.900 10.300 2.120 ;
        RECT  9.760 1.840 10.300 2.120 ;
        RECT  9.780 0.440 10.080 0.660 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.130 0.300 1.700 ;
        RECT  0.080 1.340 0.320 1.620 ;
        RECT  0.080 2.280 0.920 2.440 ;
        RECT  0.760 2.160 2.340 2.320 ;
        RECT  2.180 1.420 2.340 2.320 ;
        RECT  0.080 1.130 0.240 2.440 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 -0.280 2.360 0.400 ;
        RECT  3.870 -0.280 4.150 0.400 ;
        RECT  7.520 -0.280 7.800 0.420 ;
        RECT  9.000 -0.280 9.280 0.420 ;
        RECT  10.300 -0.280 10.580 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.320 -0.280 0.600 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 2.800 1.680 3.480 ;
        RECT  3.360 2.800 3.640 3.480 ;
        RECT  4.060 2.800 4.340 3.480 ;
        RECT  7.390 2.800 7.670 3.480 ;
        RECT  8.440 2.800 9.160 3.480 ;
        RECT  10.300 2.620 10.580 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.320 2.610 0.600 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.480 2.600 6.470 2.760 ;
        RECT  6.310 2.160 6.470 2.760 ;
        RECT  9.380 2.300 9.720 2.720 ;
        RECT  8.530 2.480 9.720 2.640 ;
        RECT  5.480 0.460 5.640 2.760 ;
        RECT  8.530 1.860 8.690 2.640 ;
        RECT  9.380 2.300 10.680 2.460 ;
        RECT  10.520 1.210 10.680 2.460 ;
        RECT  5.060 2.300 5.640 2.460 ;
        RECT  6.310 2.160 6.850 2.320 ;
        RECT  6.690 1.860 6.850 2.320 ;
        RECT  9.400 0.860 9.560 2.720 ;
        RECT  6.690 1.860 8.690 2.020 ;
        RECT  9.390 0.860 9.720 1.080 ;
        RECT  5.360 0.460 5.640 0.680 ;
        RECT  8.940 0.580 9.100 2.080 ;
        RECT  8.940 1.340 9.240 1.620 ;
        RECT  8.400 0.580 9.100 0.740 ;
        RECT  5.800 2.180 6.150 2.440 ;
        RECT  5.800 0.460 5.960 2.440 ;
        RECT  8.600 1.140 8.760 1.660 ;
        RECT  6.440 1.140 8.760 1.300 ;
        RECT  6.440 0.460 6.600 1.300 ;
        RECT  5.800 0.460 6.600 0.620 ;
        RECT  7.960 0.580 8.240 0.980 ;
        RECT  6.760 0.580 8.240 0.740 ;
        RECT  6.760 0.460 7.360 0.740 ;
        RECT  6.720 2.480 7.250 2.640 ;
        RECT  7.960 2.180 8.240 2.520 ;
        RECT  7.090 2.360 8.240 2.520 ;
        RECT  6.120 1.460 6.520 1.980 ;
        RECT  6.120 1.460 8.100 1.620 ;
        RECT  6.120 0.840 6.280 1.980 ;
        RECT  2.480 2.540 2.760 2.760 ;
        RECT  2.500 1.460 2.660 2.760 ;
        RECT  5.160 0.880 5.320 2.080 ;
        RECT  2.500 1.460 3.380 1.620 ;
        RECT  3.220 0.440 3.380 1.620 ;
        RECT  5.040 0.440 5.200 1.040 ;
        RECT  1.190 0.560 4.500 0.720 ;
        RECT  4.340 0.440 5.200 0.600 ;
        RECT  2.960 0.440 3.380 0.720 ;
        RECT  0.840 0.440 1.350 0.600 ;
        RECT  4.680 0.760 4.840 2.340 ;
        RECT  4.680 1.380 4.980 1.660 ;
        RECT  3.680 2.140 3.900 2.420 ;
        RECT  3.680 2.140 4.500 2.300 ;
        RECT  4.340 0.920 4.500 2.300 ;
        RECT  3.580 0.920 4.500 1.080 ;
        RECT  0.400 1.840 0.600 2.120 ;
        RECT  0.520 0.880 0.680 2.000 ;
        RECT  2.780 0.880 3.060 1.300 ;
        RECT  1.860 0.880 2.140 1.200 ;
        RECT  0.520 0.880 3.060 1.040 ;
        RECT  0.800 2.600 1.240 2.760 ;
        RECT  1.080 2.480 2.280 2.640 ;
    END
END DFZCRBEHD

MACRO DFZCRBHHD
    CLASS CORE ;
    FOREIGN DFZCRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.420 1.900 2.000 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.350 4.010 1.630 ;
        RECT  3.700 1.240 3.900 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.890 3.500 2.460 ;
        RECT  3.290 1.900 3.500 2.180 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 0.840 11.900 2.360 ;
        RECT  11.560 2.080 11.900 2.360 ;
        RECT  11.560 0.840 11.900 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 2.000 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.700 2.260 ;
        RECT  10.440 1.980 10.700 2.260 ;
        RECT  10.440 0.960 10.700 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.080 1.130 0.300 1.700 ;
        RECT  0.080 1.340 0.320 1.620 ;
        RECT  0.080 2.280 0.920 2.440 ;
        RECT  0.760 2.160 2.340 2.320 ;
        RECT  2.180 1.420 2.340 2.320 ;
        RECT  0.080 1.130 0.240 2.440 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 -0.280 2.360 0.400 ;
        RECT  3.870 -0.280 4.150 0.400 ;
        RECT  7.520 -0.280 7.800 0.420 ;
        RECT  8.360 -0.280 8.640 0.420 ;
        RECT  9.820 -0.280 10.100 0.400 ;
        RECT  10.940 -0.280 11.220 0.400 ;
        RECT  12.020 -0.280 12.300 0.580 ;
        RECT  0.000 -0.280 12.400 0.280 ;
        RECT  0.320 -0.280 0.600 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 2.800 1.680 3.480 ;
        RECT  3.360 2.800 3.640 3.480 ;
        RECT  4.060 2.800 4.340 3.480 ;
        RECT  7.390 2.800 7.670 3.480 ;
        RECT  8.360 2.800 8.640 3.480 ;
        RECT  9.820 2.800 10.100 3.480 ;
        RECT  10.940 2.800 11.220 3.480 ;
        RECT  12.020 2.620 12.300 3.480 ;
        RECT  0.000 2.920 12.400 3.480 ;
        RECT  0.320 2.610 0.600 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.480 2.600 6.470 2.760 ;
        RECT  6.310 2.160 6.470 2.760 ;
        RECT  8.450 2.440 11.400 2.600 ;
        RECT  11.240 0.560 11.400 2.600 ;
        RECT  5.480 0.460 5.640 2.760 ;
        RECT  5.060 2.300 5.640 2.460 ;
        RECT  8.450 1.860 8.610 2.600 ;
        RECT  6.310 2.160 6.850 2.320 ;
        RECT  6.690 1.860 6.850 2.320 ;
        RECT  6.690 1.860 8.610 2.020 ;
        RECT  9.260 0.540 9.540 0.760 ;
        RECT  9.260 0.560 11.400 0.720 ;
        RECT  5.360 0.460 5.640 0.680 ;
        RECT  8.860 1.840 9.140 2.120 ;
        RECT  8.860 0.960 9.020 2.120 ;
        RECT  8.860 1.480 9.920 1.640 ;
        RECT  8.860 0.960 9.140 1.240 ;
        RECT  5.800 2.180 6.150 2.440 ;
        RECT  5.800 0.460 5.960 2.440 ;
        RECT  8.520 1.140 8.680 1.690 ;
        RECT  6.440 1.140 8.680 1.300 ;
        RECT  6.440 0.460 6.600 1.300 ;
        RECT  5.800 0.460 6.600 0.620 ;
        RECT  7.960 0.580 8.240 0.980 ;
        RECT  6.760 0.580 8.240 0.740 ;
        RECT  6.760 0.460 7.360 0.740 ;
        RECT  6.720 2.480 7.250 2.640 ;
        RECT  7.960 2.180 8.240 2.520 ;
        RECT  7.090 2.360 8.240 2.520 ;
        RECT  6.120 1.460 6.520 1.980 ;
        RECT  6.120 1.460 8.100 1.620 ;
        RECT  6.120 0.840 6.280 1.980 ;
        RECT  2.480 2.540 2.760 2.760 ;
        RECT  2.500 1.460 2.660 2.760 ;
        RECT  5.160 0.880 5.320 2.080 ;
        RECT  2.500 1.460 3.380 1.620 ;
        RECT  3.220 0.440 3.380 1.620 ;
        RECT  5.040 0.440 5.200 1.040 ;
        RECT  1.190 0.560 4.500 0.720 ;
        RECT  4.340 0.440 5.200 0.600 ;
        RECT  2.960 0.440 3.380 0.720 ;
        RECT  0.840 0.440 1.350 0.600 ;
        RECT  4.680 0.760 4.840 2.340 ;
        RECT  4.680 1.380 4.980 1.660 ;
        RECT  3.680 2.140 3.900 2.420 ;
        RECT  3.680 2.140 4.500 2.300 ;
        RECT  4.340 0.920 4.500 2.300 ;
        RECT  3.580 0.920 4.500 1.080 ;
        RECT  0.400 1.840 0.600 2.120 ;
        RECT  0.520 0.880 0.680 2.000 ;
        RECT  2.780 0.880 3.060 1.300 ;
        RECT  1.860 0.880 2.140 1.200 ;
        RECT  0.520 0.880 3.060 1.040 ;
        RECT  0.800 2.600 1.240 2.760 ;
        RECT  1.080 2.480 2.280 2.640 ;
    END
END DFZCRBHHD

MACRO DFZECHD
    CLASS CORE ;
    FOREIGN DFZECHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 0.840 13.500 2.260 ;
        RECT  13.280 1.980 13.500 2.260 ;
        RECT  13.280 0.840 13.500 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.100 0.960 12.320 1.240 ;
        RECT  12.160 2.040 12.320 2.320 ;
        RECT  12.100 0.960 12.300 2.280 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.900 -0.280 6.180 0.400 ;
        RECT  11.260 -0.280 11.420 0.460 ;
        RECT  12.660 -0.280 12.940 0.400 ;
        RECT  0.000 -0.280 13.600 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  5.900 2.800 6.180 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  10.120 2.800 10.400 3.480 ;
        RECT  11.200 2.800 11.480 3.480 ;
        RECT  12.660 2.800 12.940 3.480 ;
        RECT  0.000 2.920 13.600 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.760 2.480 12.040 2.760 ;
        RECT  7.320 2.600 8.290 2.760 ;
        RECT  8.130 2.140 8.290 2.760 ;
        RECT  10.020 2.480 13.100 2.640 ;
        RECT  12.940 0.560 13.100 2.640 ;
        RECT  6.940 2.300 7.480 2.640 ;
        RECT  4.470 2.480 7.480 2.640 ;
        RECT  10.020 2.140 10.180 2.640 ;
        RECT  4.470 1.940 4.630 2.640 ;
        RECT  8.130 2.140 10.180 2.300 ;
        RECT  7.320 0.460 7.480 2.760 ;
        RECT  2.540 1.940 4.630 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  12.340 0.560 13.100 0.720 ;
        RECT  7.200 0.460 7.480 0.680 ;
        RECT  11.760 0.440 12.500 0.600 ;
        RECT  10.760 2.160 11.670 2.320 ;
        RECT  11.510 0.960 11.670 2.320 ;
        RECT  11.120 0.960 11.670 1.180 ;
        RECT  7.640 2.280 7.970 2.440 ;
        RECT  7.640 0.440 7.800 2.440 ;
        RECT  10.800 0.440 10.960 1.640 ;
        RECT  7.640 0.440 10.960 0.600 ;
        RECT  10.340 1.820 10.500 2.210 ;
        RECT  8.580 1.820 10.500 1.980 ;
        RECT  10.240 0.760 10.400 1.640 ;
        RECT  8.900 0.760 10.400 0.920 ;
        RECT  9.760 1.080 10.040 1.330 ;
        RECT  8.480 1.080 10.040 1.240 ;
        RECT  8.480 0.880 8.640 1.240 ;
        RECT  9.620 2.480 9.840 2.760 ;
        RECT  8.620 2.480 9.840 2.640 ;
        RECT  7.960 1.820 8.340 1.980 ;
        RECT  7.960 0.880 8.120 1.980 ;
        RECT  7.960 1.400 9.240 1.560 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.000 0.840 7.160 2.040 ;
        RECT  6.880 0.440 7.040 1.000 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.500 0.720 ;
        RECT  6.340 0.440 7.040 0.600 ;
        RECT  6.520 0.880 6.680 2.300 ;
        RECT  6.520 1.380 6.840 1.660 ;
        RECT  6.460 0.880 6.680 1.160 ;
        RECT  5.340 2.120 6.300 2.280 ;
        RECT  6.140 0.920 6.300 2.280 ;
        RECT  6.140 1.460 6.360 1.740 ;
        RECT  5.340 0.920 6.300 1.080 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.960 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZECHD

MACRO DFZEEHD
    CLASS CORE ;
    FOREIGN DFZEEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 0.840 13.500 2.260 ;
        RECT  13.280 1.980 13.500 2.260 ;
        RECT  13.280 0.840 13.500 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.100 0.960 12.320 1.240 ;
        RECT  12.160 2.040 12.320 2.320 ;
        RECT  12.100 0.960 12.300 2.280 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.900 -0.280 6.180 0.400 ;
        RECT  11.260 -0.280 11.420 0.460 ;
        RECT  12.660 -0.280 12.940 0.400 ;
        RECT  0.000 -0.280 13.600 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  5.900 2.800 6.180 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  10.120 2.800 10.400 3.480 ;
        RECT  11.200 2.800 11.480 3.480 ;
        RECT  12.660 2.800 12.940 3.480 ;
        RECT  0.000 2.920 13.600 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.760 2.480 12.040 2.760 ;
        RECT  7.320 2.600 8.290 2.760 ;
        RECT  8.130 2.140 8.290 2.760 ;
        RECT  10.020 2.480 13.100 2.640 ;
        RECT  12.940 0.560 13.100 2.640 ;
        RECT  6.940 2.300 7.480 2.640 ;
        RECT  4.470 2.480 7.480 2.640 ;
        RECT  10.020 2.140 10.180 2.640 ;
        RECT  4.470 1.940 4.630 2.640 ;
        RECT  8.130 2.140 10.180 2.300 ;
        RECT  7.320 0.460 7.480 2.760 ;
        RECT  2.540 1.940 4.630 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  12.340 0.560 13.100 0.720 ;
        RECT  7.200 0.460 7.480 0.680 ;
        RECT  11.760 0.440 12.500 0.600 ;
        RECT  10.760 2.160 11.670 2.320 ;
        RECT  11.510 0.960 11.670 2.320 ;
        RECT  11.120 0.960 11.670 1.180 ;
        RECT  7.640 2.280 7.970 2.440 ;
        RECT  7.640 0.440 7.800 2.440 ;
        RECT  10.800 0.440 10.960 1.640 ;
        RECT  7.640 0.440 10.960 0.600 ;
        RECT  10.340 1.820 10.500 2.210 ;
        RECT  8.580 1.820 10.500 1.980 ;
        RECT  10.240 0.760 10.400 1.640 ;
        RECT  8.900 0.760 10.400 0.920 ;
        RECT  9.760 1.080 10.040 1.330 ;
        RECT  8.480 1.080 10.040 1.240 ;
        RECT  8.480 0.880 8.640 1.240 ;
        RECT  9.620 2.480 9.840 2.760 ;
        RECT  8.620 2.480 9.840 2.640 ;
        RECT  7.960 1.820 8.340 1.980 ;
        RECT  7.960 0.880 8.120 1.980 ;
        RECT  7.960 1.400 9.240 1.560 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.000 0.840 7.160 2.040 ;
        RECT  6.880 0.440 7.040 1.000 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.500 0.720 ;
        RECT  6.340 0.440 7.040 0.600 ;
        RECT  6.520 0.880 6.680 2.300 ;
        RECT  6.520 1.380 6.840 1.660 ;
        RECT  6.460 0.880 6.680 1.160 ;
        RECT  5.340 2.160 6.300 2.320 ;
        RECT  6.140 0.920 6.300 2.320 ;
        RECT  6.140 1.460 6.360 1.740 ;
        RECT  5.340 0.920 6.300 1.080 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.960 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZEEHD

MACRO DFZEHD
    CLASS CORE ;
    FOREIGN DFZEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.350 3.190 1.630 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 0.580 10.300 2.120 ;
        RECT  10.080 1.840 10.300 2.120 ;
        RECT  10.080 0.580 10.300 0.860 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.300 9.100 2.120 ;
        RECT  9.060 0.440 9.260 1.500 ;
        RECT  8.980 0.440 9.260 0.660 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 3.330 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  8.180 -0.280 8.460 0.420 ;
        RECT  9.560 -0.280 9.780 0.660 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.520 3.480 ;
        RECT  6.570 2.800 6.850 3.480 ;
        RECT  7.620 2.800 8.360 3.480 ;
        RECT  9.500 2.620 9.780 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  8.580 2.300 8.920 2.720 ;
        RECT  7.710 2.480 8.920 2.640 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  7.710 1.860 7.870 2.640 ;
        RECT  8.580 2.300 9.880 2.460 ;
        RECT  9.720 1.210 9.880 2.460 ;
        RECT  4.240 2.300 4.820 2.460 ;
        RECT  5.490 2.160 6.030 2.320 ;
        RECT  5.870 1.860 6.030 2.320 ;
        RECT  8.580 0.860 8.740 2.720 ;
        RECT  5.870 1.860 7.870 2.020 ;
        RECT  8.570 0.860 8.900 1.080 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  8.120 0.580 8.280 2.080 ;
        RECT  8.120 1.340 8.420 1.620 ;
        RECT  7.580 0.580 8.280 0.740 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.780 1.140 7.940 1.660 ;
        RECT  5.620 1.140 7.940 1.300 ;
        RECT  5.620 0.460 5.780 1.300 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  7.140 0.580 7.420 0.980 ;
        RECT  5.940 0.580 7.420 0.740 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  5.900 2.480 6.430 2.640 ;
        RECT  7.140 2.180 7.420 2.520 ;
        RECT  6.270 2.360 7.420 2.520 ;
        RECT  5.300 1.460 5.700 1.980 ;
        RECT  5.300 1.460 7.280 1.620 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.660 0.560 3.680 0.720 ;
        RECT  3.520 0.440 4.380 0.600 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  3.860 0.760 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.920 3.680 2.310 ;
        RECT  2.760 0.920 3.680 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END DFZEHD

MACRO DFZEHHD
    CLASS CORE ;
    FOREIGN DFZEHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.100 0.840 14.300 2.260 ;
        RECT  13.960 1.980 14.300 2.260 ;
        RECT  13.960 0.840 14.300 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.900 0.960 13.100 2.320 ;
        RECT  12.840 2.040 13.100 2.320 ;
        RECT  12.840 0.960 13.100 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.900 -0.280 6.180 0.400 ;
        RECT  10.580 -0.280 10.800 0.500 ;
        RECT  12.220 -0.280 12.500 0.400 ;
        RECT  13.340 -0.280 13.620 0.400 ;
        RECT  14.420 -0.280 14.700 0.580 ;
        RECT  0.000 -0.280 14.800 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  5.900 2.800 6.180 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  11.320 2.800 11.600 3.480 ;
        RECT  12.220 2.800 12.500 3.480 ;
        RECT  13.340 2.800 13.620 3.480 ;
        RECT  14.420 2.620 14.700 3.480 ;
        RECT  0.000 2.920 14.800 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.320 2.600 8.290 2.760 ;
        RECT  8.130 2.140 8.290 2.760 ;
        RECT  10.020 2.480 13.780 2.640 ;
        RECT  13.620 0.560 13.780 2.640 ;
        RECT  6.940 2.300 7.480 2.640 ;
        RECT  4.470 2.480 7.480 2.640 ;
        RECT  11.880 2.280 12.160 2.640 ;
        RECT  10.020 2.140 10.180 2.640 ;
        RECT  4.470 1.940 4.630 2.640 ;
        RECT  8.130 2.140 10.180 2.300 ;
        RECT  7.320 0.460 7.480 2.760 ;
        RECT  2.540 1.940 4.630 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  11.660 0.560 13.780 0.720 ;
        RECT  7.200 0.460 7.480 0.680 ;
        RECT  10.760 2.160 11.670 2.320 ;
        RECT  11.510 0.960 11.670 2.320 ;
        RECT  11.080 0.960 11.670 1.180 ;
        RECT  7.640 2.280 7.970 2.440 ;
        RECT  7.640 0.440 7.800 2.440 ;
        RECT  10.780 1.270 10.940 1.680 ;
        RECT  10.260 1.270 10.940 1.430 ;
        RECT  10.260 0.440 10.420 1.430 ;
        RECT  7.640 0.440 10.420 0.600 ;
        RECT  10.340 1.820 10.500 2.210 ;
        RECT  8.580 1.820 10.500 1.980 ;
        RECT  9.940 0.760 10.100 1.660 ;
        RECT  8.900 0.760 10.100 0.920 ;
        RECT  9.620 2.480 9.840 2.760 ;
        RECT  8.620 2.480 9.840 2.640 ;
        RECT  9.500 1.080 9.780 1.330 ;
        RECT  8.480 1.080 9.780 1.240 ;
        RECT  8.480 0.880 8.640 1.240 ;
        RECT  7.960 1.820 8.340 1.980 ;
        RECT  7.960 0.880 8.120 1.980 ;
        RECT  7.960 1.400 9.240 1.560 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.000 0.840 7.160 2.040 ;
        RECT  6.880 0.440 7.040 1.000 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.500 0.720 ;
        RECT  6.340 0.440 7.040 0.600 ;
        RECT  6.520 0.880 6.680 2.300 ;
        RECT  6.520 1.380 6.840 1.660 ;
        RECT  6.460 0.880 6.680 1.160 ;
        RECT  5.340 2.160 6.300 2.320 ;
        RECT  6.140 0.920 6.300 2.320 ;
        RECT  6.140 1.460 6.360 1.740 ;
        RECT  5.340 0.920 6.300 1.080 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.960 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZEHHD

MACRO DFZEKHD
    CLASS CORE ;
    FOREIGN DFZEKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.920 0.860 16.120 1.140 ;
        RECT  14.920 2.060 16.120 2.340 ;
        RECT  15.250 0.860 15.550 2.340 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.840 0.860 14.040 1.140 ;
        RECT  12.840 1.840 14.040 2.120 ;
        RECT  13.250 0.860 13.550 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.840 -0.280 5.120 0.400 ;
        RECT  5.880 -0.280 6.160 0.400 ;
        RECT  10.560 -0.280 10.780 0.640 ;
        RECT  12.260 -0.280 12.540 0.580 ;
        RECT  13.300 -0.280 13.580 0.580 ;
        RECT  14.340 -0.280 14.620 0.580 ;
        RECT  15.380 -0.280 15.660 0.580 ;
        RECT  16.420 -0.280 16.700 0.580 ;
        RECT  0.000 -0.280 16.800 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.810 2.800 5.090 3.480 ;
        RECT  5.880 2.800 6.160 3.480 ;
        RECT  9.160 2.800 9.440 3.480 ;
        RECT  11.320 2.800 11.600 3.480 ;
        RECT  12.220 2.800 12.500 3.480 ;
        RECT  13.300 2.620 13.580 3.480 ;
        RECT  14.340 2.620 14.620 3.480 ;
        RECT  15.380 2.620 15.660 3.480 ;
        RECT  16.420 2.620 16.700 3.480 ;
        RECT  0.000 2.920 16.800 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.300 2.600 8.270 2.760 ;
        RECT  8.110 2.140 8.270 2.760 ;
        RECT  10.000 2.480 12.680 2.640 ;
        RECT  12.520 0.740 12.680 2.640 ;
        RECT  6.920 2.300 7.460 2.640 ;
        RECT  4.420 2.480 7.460 2.640 ;
        RECT  11.880 2.280 12.160 2.640 ;
        RECT  10.000 2.140 10.160 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  12.520 2.300 14.740 2.460 ;
        RECT  14.580 1.300 14.740 2.460 ;
        RECT  8.110 2.140 10.160 2.300 ;
        RECT  7.300 0.460 7.460 2.760 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  11.740 0.740 12.680 0.900 ;
        RECT  7.180 0.460 7.460 0.680 ;
        RECT  10.740 2.160 11.460 2.320 ;
        RECT  11.300 0.960 11.460 2.320 ;
        RECT  11.300 1.420 12.340 1.700 ;
        RECT  11.020 0.960 11.460 1.180 ;
        RECT  7.620 2.280 7.950 2.440 ;
        RECT  7.620 0.440 7.780 2.440 ;
        RECT  10.720 1.270 10.880 1.680 ;
        RECT  10.240 1.270 10.880 1.430 ;
        RECT  10.240 0.440 10.400 1.430 ;
        RECT  7.620 0.440 10.400 0.600 ;
        RECT  10.320 1.820 10.480 2.210 ;
        RECT  8.560 1.820 10.480 1.980 ;
        RECT  9.920 0.760 10.080 1.660 ;
        RECT  8.880 0.760 10.080 0.920 ;
        RECT  9.600 2.480 9.820 2.760 ;
        RECT  8.600 2.480 9.820 2.640 ;
        RECT  9.480 1.080 9.760 1.330 ;
        RECT  8.460 1.080 9.760 1.240 ;
        RECT  8.460 0.880 8.620 1.240 ;
        RECT  7.940 1.820 8.320 1.980 ;
        RECT  7.940 0.880 8.100 1.980 ;
        RECT  7.940 1.400 9.220 1.560 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  6.980 0.840 7.140 2.040 ;
        RECT  6.860 0.440 7.020 1.000 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.480 0.720 ;
        RECT  6.320 0.440 7.020 0.600 ;
        RECT  6.500 0.880 6.660 2.300 ;
        RECT  6.500 1.380 6.820 1.660 ;
        RECT  6.440 0.880 6.660 1.160 ;
        RECT  5.320 2.160 6.280 2.320 ;
        RECT  6.120 0.920 6.280 2.320 ;
        RECT  6.120 1.460 6.340 1.740 ;
        RECT  5.320 0.920 6.280 1.080 ;
        RECT  4.900 0.880 5.060 2.320 ;
        RECT  2.960 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.120 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZEKHD

MACRO DFZERBCHD
    CLASS CORE ;
    FOREIGN DFZERBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.200 10.890 1.660 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.680 1.840 13.900 2.120 ;
        RECT  13.700 0.920 13.900 2.160 ;
        RECT  13.680 0.960 13.900 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 0.980 12.860 2.060 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.860 -0.280 6.140 0.400 ;
        RECT  9.700 -0.280 9.980 0.400 ;
        RECT  10.780 -0.280 11.060 0.400 ;
        RECT  11.620 -0.280 11.900 0.400 ;
        RECT  13.100 -0.280 13.380 0.940 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  9.480 2.800 9.760 3.480 ;
        RECT  10.300 2.800 10.580 3.480 ;
        RECT  11.420 2.800 11.700 3.480 ;
        RECT  13.060 2.620 13.340 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.440 2.600 8.670 2.760 ;
        RECT  8.510 2.160 8.670 2.760 ;
        RECT  7.060 2.300 7.600 2.640 ;
        RECT  4.420 2.480 7.600 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  12.180 2.220 13.430 2.380 ;
        RECT  13.270 1.290 13.430 2.380 ;
        RECT  8.510 2.160 12.340 2.320 ;
        RECT  7.440 0.460 7.600 2.760 ;
        RECT  12.180 0.440 12.340 2.380 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  13.270 1.340 13.480 1.620 ;
        RECT  7.280 0.460 7.600 0.680 ;
        RECT  12.180 0.440 12.500 0.600 ;
        RECT  11.860 2.600 12.200 2.760 ;
        RECT  10.820 2.480 12.020 2.640 ;
        RECT  11.860 0.880 12.020 1.760 ;
        RECT  11.600 0.880 12.020 1.160 ;
        RECT  8.070 2.280 8.350 2.440 ;
        RECT  8.110 1.840 8.270 2.440 ;
        RECT  8.110 1.840 9.000 2.000 ;
        RECT  8.840 1.060 9.000 2.000 ;
        RECT  11.340 1.350 11.500 1.900 ;
        RECT  8.840 1.500 10.340 1.660 ;
        RECT  10.180 0.880 10.340 1.660 ;
        RECT  11.270 0.880 11.430 1.510 ;
        RECT  8.420 1.060 9.000 1.220 ;
        RECT  8.420 0.600 8.580 1.220 ;
        RECT  10.180 0.880 11.430 1.040 ;
        RECT  7.800 0.600 8.580 0.760 ;
        RECT  7.800 0.460 8.140 0.760 ;
        RECT  9.160 1.820 11.180 1.980 ;
        RECT  9.240 0.560 10.400 0.720 ;
        RECT  10.140 0.440 10.400 0.720 ;
        RECT  8.770 0.460 9.400 0.620 ;
        RECT  8.830 2.480 10.190 2.640 ;
        RECT  9.160 0.880 10.020 1.160 ;
        RECT  7.760 0.940 7.920 2.080 ;
        RECT  7.760 1.380 8.680 1.660 ;
        RECT  7.760 0.940 8.120 1.100 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.120 0.880 7.280 2.080 ;
        RECT  6.960 0.440 7.120 1.040 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.460 0.720 ;
        RECT  6.300 0.440 7.120 0.600 ;
        RECT  6.640 0.760 6.800 2.320 ;
        RECT  6.640 1.380 6.940 1.660 ;
        RECT  5.540 2.160 6.460 2.320 ;
        RECT  6.300 0.880 6.460 2.320 ;
        RECT  5.540 0.880 6.460 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERBCHD

MACRO DFZERBEHD
    CLASS CORE ;
    FOREIGN DFZERBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 1.200 10.540 1.660 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 1.420 5.600 1.700 ;
        RECT  5.300 1.420 5.500 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.680 1.840 13.900 2.120 ;
        RECT  13.700 0.920 13.900 2.160 ;
        RECT  13.680 0.960 13.900 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 1.840 12.780 2.120 ;
        RECT  12.500 1.020 12.860 1.240 ;
        RECT  12.500 0.980 12.700 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.800 -0.280 5.080 0.400 ;
        RECT  5.560 -0.280 5.840 0.400 ;
        RECT  9.400 -0.280 9.680 0.400 ;
        RECT  10.480 -0.280 10.760 0.400 ;
        RECT  11.700 -0.280 11.980 0.580 ;
        RECT  13.100 -0.280 13.380 0.580 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.770 2.800 5.050 3.480 ;
        RECT  5.720 2.800 6.000 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  10.000 2.800 10.280 3.480 ;
        RECT  11.160 2.800 11.440 3.480 ;
        RECT  13.100 2.620 13.380 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.140 2.600 8.370 2.760 ;
        RECT  8.210 2.160 8.370 2.760 ;
        RECT  6.760 2.300 7.300 2.640 ;
        RECT  4.420 2.480 7.300 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  12.160 2.300 13.430 2.460 ;
        RECT  13.270 1.340 13.430 2.460 ;
        RECT  8.210 2.160 12.320 2.320 ;
        RECT  7.140 0.460 7.300 2.760 ;
        RECT  12.160 0.440 12.320 2.460 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  13.270 1.340 13.480 1.620 ;
        RECT  12.160 0.440 12.500 0.750 ;
        RECT  6.980 0.460 7.300 0.680 ;
        RECT  11.840 0.880 12.000 1.480 ;
        RECT  11.420 0.880 12.000 1.160 ;
        RECT  11.600 2.480 11.880 2.740 ;
        RECT  10.520 2.480 11.880 2.640 ;
        RECT  7.770 2.280 8.050 2.440 ;
        RECT  7.810 1.840 7.970 2.440 ;
        RECT  7.810 1.840 8.700 2.000 ;
        RECT  8.540 1.060 8.700 2.000 ;
        RECT  11.100 1.440 11.520 1.720 ;
        RECT  8.540 1.500 9.940 1.660 ;
        RECT  9.780 0.880 9.940 1.660 ;
        RECT  11.100 0.880 11.260 1.720 ;
        RECT  8.120 1.060 8.700 1.220 ;
        RECT  8.120 0.600 8.280 1.220 ;
        RECT  9.780 0.880 11.260 1.040 ;
        RECT  7.500 0.600 8.280 0.760 ;
        RECT  7.500 0.460 7.840 0.760 ;
        RECT  8.860 1.820 10.880 1.980 ;
        RECT  8.940 0.560 10.100 0.720 ;
        RECT  9.840 0.440 10.100 0.720 ;
        RECT  8.470 0.460 9.100 0.620 ;
        RECT  8.530 2.480 9.890 2.640 ;
        RECT  8.860 0.880 9.620 1.160 ;
        RECT  7.460 0.940 7.620 2.080 ;
        RECT  7.460 1.380 8.380 1.660 ;
        RECT  7.460 0.940 7.820 1.100 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  6.820 0.880 6.980 2.080 ;
        RECT  6.660 0.440 6.820 1.040 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.160 0.720 ;
        RECT  6.000 0.440 6.820 0.600 ;
        RECT  6.340 0.760 6.500 2.320 ;
        RECT  6.340 1.380 6.640 1.660 ;
        RECT  5.200 2.160 6.160 2.320 ;
        RECT  6.000 0.880 6.160 2.320 ;
        RECT  5.240 0.880 6.160 1.040 ;
        RECT  4.860 0.880 5.020 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.020 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERBEHD

MACRO DFZERBHHD
    CLASS CORE ;
    FOREIGN DFZERBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.200 10.890 1.660 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.900 0.920 15.100 2.160 ;
        RECT  14.720 1.840 15.100 2.160 ;
        RECT  14.720 0.920 15.100 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.700 0.960 13.900 2.120 ;
        RECT  13.680 1.840 13.900 2.120 ;
        RECT  13.680 0.960 13.900 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.860 -0.280 6.140 0.400 ;
        RECT  9.700 -0.280 9.980 0.400 ;
        RECT  10.780 -0.280 11.440 0.580 ;
        RECT  13.100 -0.280 13.380 0.580 ;
        RECT  14.140 -0.280 14.420 0.580 ;
        RECT  15.180 -0.280 15.460 0.580 ;
        RECT  0.000 -0.280 15.600 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  9.480 2.800 9.760 3.480 ;
        RECT  10.280 2.800 10.560 3.480 ;
        RECT  11.200 2.620 11.480 3.480 ;
        RECT  12.240 2.620 12.520 3.480 ;
        RECT  13.100 2.620 13.380 3.480 ;
        RECT  14.140 2.620 14.420 3.480 ;
        RECT  15.180 2.620 15.460 3.480 ;
        RECT  0.000 2.920 15.600 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.440 2.600 8.670 2.760 ;
        RECT  8.510 2.160 8.670 2.760 ;
        RECT  7.060 2.300 7.600 2.640 ;
        RECT  4.430 2.480 7.600 2.640 ;
        RECT  4.430 1.940 4.590 2.640 ;
        RECT  10.370 2.300 14.470 2.460 ;
        RECT  14.310 1.340 14.470 2.460 ;
        RECT  8.510 2.160 10.530 2.320 ;
        RECT  12.640 2.020 12.920 2.460 ;
        RECT  12.760 0.780 12.920 2.460 ;
        RECT  7.440 0.460 7.600 2.760 ;
        RECT  2.540 1.940 4.590 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  14.310 1.340 14.520 1.620 ;
        RECT  12.640 0.780 12.920 1.060 ;
        RECT  7.280 0.460 7.600 0.680 ;
        RECT  11.680 1.950 12.480 2.110 ;
        RECT  12.320 0.490 12.480 2.110 ;
        RECT  12.320 1.460 12.600 1.740 ;
        RECT  12.000 0.490 12.480 0.650 ;
        RECT  8.070 2.280 8.350 2.440 ;
        RECT  8.110 1.840 8.270 2.440 ;
        RECT  8.110 1.840 9.000 2.000 ;
        RECT  8.840 1.060 9.000 2.000 ;
        RECT  11.960 0.880 12.120 1.670 ;
        RECT  8.840 1.500 10.340 1.660 ;
        RECT  10.180 0.880 10.340 1.660 ;
        RECT  8.420 1.060 9.000 1.220 ;
        RECT  8.420 0.600 8.580 1.220 ;
        RECT  10.180 0.880 12.120 1.040 ;
        RECT  7.800 0.600 8.580 0.760 ;
        RECT  7.800 0.460 8.140 0.760 ;
        RECT  10.860 1.820 11.140 2.140 ;
        RECT  9.160 1.820 11.140 1.980 ;
        RECT  9.240 0.560 10.400 0.720 ;
        RECT  10.140 0.440 10.400 0.720 ;
        RECT  8.770 0.460 9.400 0.620 ;
        RECT  8.830 2.480 10.190 2.640 ;
        RECT  9.160 0.880 10.020 1.160 ;
        RECT  7.760 0.940 7.920 2.080 ;
        RECT  7.760 1.380 8.680 1.660 ;
        RECT  7.760 0.940 8.120 1.100 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.120 0.880 7.280 2.080 ;
        RECT  6.960 0.440 7.120 1.040 ;
        RECT  1.600 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.460 0.720 ;
        RECT  6.300 0.440 7.120 0.600 ;
        RECT  6.640 0.760 6.800 2.320 ;
        RECT  6.640 1.380 6.940 1.660 ;
        RECT  5.540 2.160 6.460 2.320 ;
        RECT  6.300 0.880 6.460 2.320 ;
        RECT  5.540 0.880 6.460 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERBHHD

MACRO DFZERBKHD
    CLASS CORE ;
    FOREIGN DFZERBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 1.200 11.500 1.960 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.200 5.900 1.800 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.720 0.960 16.920 1.240 ;
        RECT  15.720 1.840 16.920 2.120 ;
        RECT  16.050 0.960 16.350 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.640 0.960 14.840 1.240 ;
        RECT  13.640 1.840 14.840 2.120 ;
        RECT  14.050 0.960 14.350 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.720 -0.280 5.000 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  10.370 -0.280 10.970 0.460 ;
        RECT  11.190 -0.280 11.470 0.580 ;
        RECT  13.060 -0.280 13.340 0.580 ;
        RECT  14.100 -0.280 14.380 0.580 ;
        RECT  15.140 -0.280 15.420 0.580 ;
        RECT  16.180 -0.280 16.460 0.580 ;
        RECT  17.220 -0.280 17.500 0.580 ;
        RECT  0.000 -0.280 17.600 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.870 2.800 5.150 3.480 ;
        RECT  6.140 2.800 6.420 3.480 ;
        RECT  9.260 2.800 9.540 3.480 ;
        RECT  10.360 2.800 10.640 3.480 ;
        RECT  11.120 2.800 11.400 3.480 ;
        RECT  12.200 2.620 12.480 3.480 ;
        RECT  13.060 2.620 13.340 3.480 ;
        RECT  14.100 2.620 14.380 3.480 ;
        RECT  15.140 2.620 15.420 3.480 ;
        RECT  16.180 2.620 16.460 3.480 ;
        RECT  17.220 2.620 17.500 3.480 ;
        RECT  0.000 2.920 17.600 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 2.600 8.530 2.760 ;
        RECT  8.370 2.160 8.530 2.760 ;
        RECT  7.180 2.300 7.720 2.640 ;
        RECT  4.420 2.480 7.720 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  10.490 2.300 15.470 2.460 ;
        RECT  15.310 1.340 15.470 2.460 ;
        RECT  8.370 2.160 10.650 2.320 ;
        RECT  12.600 2.020 12.880 2.460 ;
        RECT  12.720 0.960 12.880 2.460 ;
        RECT  7.560 0.460 7.720 2.760 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  15.310 1.340 15.520 1.620 ;
        RECT  12.600 0.960 12.880 1.240 ;
        RECT  7.400 0.460 7.720 0.680 ;
        RECT  11.680 1.950 12.440 2.110 ;
        RECT  12.280 0.490 12.440 2.110 ;
        RECT  11.680 1.890 11.960 2.110 ;
        RECT  12.280 1.460 12.560 1.740 ;
        RECT  11.990 0.490 12.440 0.650 ;
        RECT  7.880 2.220 8.210 2.440 ;
        RECT  7.880 0.440 8.040 2.440 ;
        RECT  11.910 0.810 12.070 1.670 ;
        RECT  10.740 0.810 12.070 0.970 ;
        RECT  10.740 0.620 10.900 0.970 ;
        RECT  10.050 0.620 10.900 0.780 ;
        RECT  10.050 0.440 10.210 0.780 ;
        RECT  7.880 0.440 10.210 0.600 ;
        RECT  10.820 1.820 11.100 2.140 ;
        RECT  8.780 1.820 11.100 1.980 ;
        RECT  9.410 1.380 10.440 1.540 ;
        RECT  10.280 0.940 10.440 1.540 ;
        RECT  9.410 1.120 9.570 1.540 ;
        RECT  8.660 1.120 9.570 1.280 ;
        RECT  10.280 0.940 10.560 1.160 ;
        RECT  8.660 0.940 8.940 1.280 ;
        RECT  8.700 2.480 8.980 2.700 ;
        RECT  8.700 2.480 10.300 2.640 ;
        RECT  9.730 0.940 10.060 1.220 ;
        RECT  9.730 0.760 9.890 1.220 ;
        RECT  9.100 0.760 9.890 0.920 ;
        RECT  8.200 1.440 8.580 1.980 ;
        RECT  8.970 1.440 9.250 1.660 ;
        RECT  8.200 1.440 9.250 1.600 ;
        RECT  8.200 0.840 8.360 1.980 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.240 0.880 7.400 2.080 ;
        RECT  7.080 0.560 7.240 1.040 ;
        RECT  1.590 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 7.240 0.720 ;
        RECT  6.760 0.880 6.920 2.320 ;
        RECT  6.760 1.380 7.060 1.660 ;
        RECT  6.700 0.880 6.920 1.160 ;
        RECT  5.540 2.160 6.540 2.320 ;
        RECT  6.380 0.880 6.540 2.320 ;
        RECT  6.380 1.460 6.580 1.740 ;
        RECT  5.540 0.880 6.540 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.080 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERBKHD

MACRO DFZERSBCHD
    CLASS CORE ;
    FOREIGN DFZERSBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.090 0.840 11.500 1.340 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.880 1.840 15.100 2.120 ;
        RECT  14.900 0.920 15.100 2.160 ;
        RECT  14.880 0.960 15.100 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.700 1.840 13.920 2.120 ;
        RECT  13.700 1.020 14.060 1.240 ;
        RECT  13.700 0.980 13.900 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 1.380 12.700 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.860 -0.280 6.140 0.400 ;
        RECT  9.980 -0.280 10.260 0.620 ;
        RECT  11.380 -0.280 11.660 0.620 ;
        RECT  12.600 -0.280 12.880 0.620 ;
        RECT  14.300 -0.280 14.580 0.940 ;
        RECT  0.000 -0.280 15.200 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  9.480 2.800 9.760 3.480 ;
        RECT  10.960 2.800 11.240 3.480 ;
        RECT  12.200 2.800 12.480 3.480 ;
        RECT  13.220 2.800 13.500 3.480 ;
        RECT  14.260 2.620 14.540 3.480 ;
        RECT  0.000 2.920 15.200 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.440 2.600 8.670 2.760 ;
        RECT  8.510 2.160 8.670 2.760 ;
        RECT  7.060 2.300 7.600 2.640 ;
        RECT  4.420 2.480 7.600 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  13.380 2.300 14.630 2.460 ;
        RECT  14.470 1.340 14.630 2.460 ;
        RECT  8.510 2.160 13.540 2.320 ;
        RECT  7.440 0.460 7.600 2.760 ;
        RECT  13.380 0.440 13.540 2.460 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  14.470 1.340 14.680 1.620 ;
        RECT  13.380 0.440 13.720 0.750 ;
        RECT  7.280 0.460 7.600 0.680 ;
        RECT  13.060 0.940 13.220 1.480 ;
        RECT  12.220 0.940 13.220 1.100 ;
        RECT  12.730 2.480 13.060 2.740 ;
        RECT  11.560 2.480 13.060 2.640 ;
        RECT  8.070 2.280 8.350 2.440 ;
        RECT  8.110 1.840 8.270 2.440 ;
        RECT  8.110 1.840 9.000 2.000 ;
        RECT  8.840 1.060 9.000 2.000 ;
        RECT  12.000 1.500 12.160 1.920 ;
        RECT  8.840 1.500 12.160 1.660 ;
        RECT  8.420 1.060 9.000 1.220 ;
        RECT  8.420 0.600 8.580 1.220 ;
        RECT  7.800 0.600 8.580 0.760 ;
        RECT  7.800 0.460 8.140 0.760 ;
        RECT  9.160 1.820 11.840 1.980 ;
        RECT  8.830 2.480 10.780 2.640 ;
        RECT  9.270 1.180 10.720 1.340 ;
        RECT  10.560 0.700 10.720 1.340 ;
        RECT  9.270 0.880 9.430 1.340 ;
        RECT  9.160 0.880 9.430 1.160 ;
        RECT  9.590 0.780 10.400 1.000 ;
        RECT  9.590 0.460 9.750 1.000 ;
        RECT  8.770 0.460 9.750 0.620 ;
        RECT  7.760 0.940 7.920 2.080 ;
        RECT  7.760 1.380 8.680 1.660 ;
        RECT  7.760 0.940 8.120 1.100 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.120 0.880 7.280 2.080 ;
        RECT  6.960 0.440 7.120 1.040 ;
        RECT  1.590 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.460 0.720 ;
        RECT  6.300 0.440 7.120 0.600 ;
        RECT  6.640 0.760 6.800 2.320 ;
        RECT  6.640 1.380 6.940 1.660 ;
        RECT  5.540 2.150 6.460 2.310 ;
        RECT  6.300 0.880 6.460 2.310 ;
        RECT  5.540 0.880 6.460 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERSBCHD

MACRO DFZERSBEHD
    CLASS CORE ;
    FOREIGN DFZERSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.090 0.840 11.500 1.340 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.880 1.840 15.100 2.120 ;
        RECT  14.900 0.920 15.100 2.160 ;
        RECT  14.880 0.960 15.100 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.700 1.840 13.980 2.120 ;
        RECT  13.700 1.020 14.060 1.240 ;
        RECT  13.700 0.980 13.900 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 1.380 12.700 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.860 -0.280 6.140 0.400 ;
        RECT  9.980 -0.280 10.260 0.620 ;
        RECT  11.380 -0.280 11.660 0.620 ;
        RECT  12.600 -0.280 12.880 0.620 ;
        RECT  14.300 -0.280 14.580 0.580 ;
        RECT  0.000 -0.280 15.200 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  9.480 2.800 9.760 3.480 ;
        RECT  10.960 2.800 11.240 3.480 ;
        RECT  12.200 2.800 12.480 3.480 ;
        RECT  13.220 2.800 13.500 3.480 ;
        RECT  14.300 2.620 14.580 3.480 ;
        RECT  0.000 2.920 15.200 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.440 2.600 8.670 2.760 ;
        RECT  8.510 2.160 8.670 2.760 ;
        RECT  7.060 2.300 7.600 2.640 ;
        RECT  4.520 2.480 7.600 2.640 ;
        RECT  4.520 1.940 4.680 2.640 ;
        RECT  13.380 2.300 14.630 2.460 ;
        RECT  14.470 1.340 14.630 2.460 ;
        RECT  8.510 2.160 13.540 2.320 ;
        RECT  7.440 0.460 7.600 2.760 ;
        RECT  13.380 0.440 13.540 2.460 ;
        RECT  2.540 1.940 4.680 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  14.470 1.340 14.680 1.620 ;
        RECT  13.380 0.440 13.720 0.750 ;
        RECT  7.280 0.460 7.600 0.680 ;
        RECT  13.060 0.940 13.220 1.480 ;
        RECT  12.220 0.940 13.220 1.100 ;
        RECT  12.730 2.480 13.060 2.740 ;
        RECT  11.560 2.480 13.060 2.640 ;
        RECT  8.070 2.280 8.350 2.440 ;
        RECT  8.110 1.840 8.270 2.440 ;
        RECT  8.110 1.840 9.000 2.000 ;
        RECT  8.840 1.060 9.000 2.000 ;
        RECT  12.000 1.500 12.160 1.920 ;
        RECT  8.840 1.500 12.160 1.660 ;
        RECT  8.420 1.060 9.000 1.220 ;
        RECT  8.420 0.600 8.580 1.220 ;
        RECT  7.800 0.600 8.580 0.760 ;
        RECT  7.800 0.460 8.140 0.760 ;
        RECT  9.160 1.820 11.840 1.980 ;
        RECT  8.830 2.480 10.780 2.640 ;
        RECT  9.270 1.180 10.720 1.340 ;
        RECT  10.560 0.700 10.720 1.340 ;
        RECT  9.270 0.880 9.430 1.340 ;
        RECT  9.160 0.880 9.430 1.160 ;
        RECT  9.590 0.780 10.400 1.000 ;
        RECT  9.590 0.460 9.750 1.000 ;
        RECT  8.770 0.460 9.750 0.620 ;
        RECT  7.760 0.940 7.920 2.080 ;
        RECT  7.760 1.380 8.680 1.660 ;
        RECT  7.760 0.940 8.120 1.100 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.120 0.880 7.280 2.080 ;
        RECT  6.960 0.440 7.120 1.040 ;
        RECT  1.590 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.460 0.720 ;
        RECT  6.300 0.440 7.120 0.600 ;
        RECT  6.640 0.760 6.800 2.320 ;
        RECT  6.640 1.380 6.940 1.660 ;
        RECT  5.540 2.160 6.460 2.320 ;
        RECT  6.300 0.880 6.460 2.320 ;
        RECT  5.540 0.880 6.460 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERSBEHD

MACRO DFZERSBHHD
    CLASS CORE ;
    FOREIGN DFZERSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 1.620 11.920 1.900 ;
        RECT  11.700 1.440 11.900 1.940 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.100 0.920 16.300 2.160 ;
        RECT  15.960 1.840 16.300 2.160 ;
        RECT  15.960 0.920 16.300 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.860 0.960 15.140 1.240 ;
        RECT  14.860 1.840 15.140 2.120 ;
        RECT  14.900 0.960 15.100 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 1.420 13.500 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.860 -0.280 5.140 0.400 ;
        RECT  5.860 -0.280 6.140 0.400 ;
        RECT  10.030 -0.280 10.250 0.680 ;
        RECT  11.800 -0.280 12.080 0.620 ;
        RECT  13.120 -0.280 13.400 0.620 ;
        RECT  14.300 -0.280 14.580 0.400 ;
        RECT  15.380 -0.280 15.660 0.580 ;
        RECT  16.420 -0.280 16.700 0.580 ;
        RECT  0.000 -0.280 16.800 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.830 2.800 5.110 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  9.480 2.800 9.760 3.480 ;
        RECT  11.100 2.800 11.380 3.480 ;
        RECT  11.980 2.800 12.260 3.480 ;
        RECT  13.180 2.800 13.460 3.480 ;
        RECT  14.300 2.800 14.580 3.480 ;
        RECT  15.380 2.620 15.660 3.480 ;
        RECT  16.420 2.620 16.700 3.480 ;
        RECT  0.000 2.920 16.800 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.440 2.600 8.670 2.760 ;
        RECT  8.510 2.160 8.670 2.760 ;
        RECT  11.010 2.480 15.150 2.640 ;
        RECT  14.990 2.280 15.150 2.640 ;
        RECT  7.060 2.300 7.600 2.640 ;
        RECT  4.420 2.480 7.600 2.640 ;
        RECT  14.520 0.900 14.680 2.640 ;
        RECT  11.010 2.160 11.170 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  14.990 2.280 15.800 2.440 ;
        RECT  15.640 1.300 15.800 2.440 ;
        RECT  8.510 2.160 11.170 2.320 ;
        RECT  7.440 0.460 7.600 2.760 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  14.020 0.900 14.680 1.060 ;
        RECT  14.020 0.750 14.240 1.060 ;
        RECT  7.280 0.460 7.600 0.680 ;
        RECT  12.540 2.160 14.280 2.320 ;
        RECT  14.120 1.240 14.280 2.320 ;
        RECT  13.680 1.240 14.280 1.400 ;
        RECT  13.680 0.780 13.840 1.400 ;
        RECT  12.640 0.780 12.960 1.040 ;
        RECT  12.640 0.780 13.840 0.940 ;
        RECT  8.070 2.280 8.350 2.440 ;
        RECT  8.110 1.840 8.270 2.440 ;
        RECT  8.110 1.840 9.000 2.000 ;
        RECT  8.840 1.060 9.000 2.000 ;
        RECT  12.860 1.200 13.020 1.940 ;
        RECT  8.840 1.500 11.520 1.660 ;
        RECT  11.360 0.880 11.520 1.660 ;
        RECT  12.280 1.200 13.020 1.360 ;
        RECT  8.420 1.060 9.000 1.220 ;
        RECT  12.280 0.880 12.440 1.360 ;
        RECT  8.420 0.600 8.580 1.220 ;
        RECT  11.360 0.880 12.440 1.040 ;
        RECT  7.800 0.600 8.580 0.760 ;
        RECT  7.800 0.460 8.140 0.760 ;
        RECT  11.330 2.160 11.950 2.320 ;
        RECT  11.330 1.820 11.490 2.320 ;
        RECT  9.160 1.820 11.490 1.980 ;
        RECT  9.590 0.840 10.660 1.000 ;
        RECT  10.500 0.560 10.660 1.000 ;
        RECT  9.590 0.460 9.750 1.000 ;
        RECT  10.500 0.560 11.380 0.720 ;
        RECT  8.770 0.460 9.750 0.620 ;
        RECT  9.270 1.180 11.200 1.340 ;
        RECT  10.950 0.880 11.200 1.340 ;
        RECT  9.270 0.880 9.430 1.340 ;
        RECT  9.160 0.880 9.430 1.160 ;
        RECT  8.830 2.480 10.850 2.640 ;
        RECT  7.760 0.940 7.920 2.080 ;
        RECT  7.760 1.380 8.680 1.660 ;
        RECT  7.760 0.940 8.120 1.100 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.120 0.880 7.280 2.040 ;
        RECT  6.960 0.440 7.120 1.040 ;
        RECT  1.580 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 6.460 0.720 ;
        RECT  6.300 0.440 7.120 0.600 ;
        RECT  6.640 0.760 6.800 2.320 ;
        RECT  6.640 1.380 6.940 1.660 ;
        RECT  5.540 2.160 6.460 2.320 ;
        RECT  6.300 0.880 6.460 2.320 ;
        RECT  5.540 0.880 6.460 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.140 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERSBHHD

MACRO DFZERSBKHD
    CLASS CORE ;
    FOREIGN DFZERSBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 1.350 11.900 1.940 ;
        RECT  11.680 1.620 11.900 1.900 ;
        END
    END RB
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.300 0.300 1.960 ;
        END
    END EB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.420 5.970 1.700 ;
        RECT  5.700 1.420 5.900 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.200 4.300 1.740 ;
        RECT  4.060 1.420 4.300 1.700 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  16.920 0.960 18.120 1.240 ;
        RECT  16.920 1.840 18.120 2.120 ;
        RECT  17.250 0.960 17.550 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.140 1.580 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.840 0.960 16.040 1.240 ;
        RECT  14.840 1.840 16.040 2.120 ;
        RECT  15.250 0.960 15.550 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 1.260 13.500 1.960 ;
        RECT  13.280 1.420 13.500 1.700 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.200 4.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.400 ;
        RECT  4.720 -0.280 5.000 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  10.060 -0.280 10.340 0.400 ;
        RECT  11.720 -0.280 12.000 0.620 ;
        RECT  13.040 -0.280 13.320 0.620 ;
        RECT  14.220 -0.280 14.500 0.400 ;
        RECT  15.300 -0.280 15.580 0.580 ;
        RECT  16.340 -0.280 16.620 0.580 ;
        RECT  17.380 -0.280 17.660 0.580 ;
        RECT  18.420 -0.280 18.700 0.580 ;
        RECT  0.000 -0.280 18.800 0.280 ;
        RECT  0.320 -0.280 0.600 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 2.580 3.380 3.480 ;
        RECT  4.870 2.800 5.150 3.480 ;
        RECT  6.140 2.800 6.420 3.480 ;
        RECT  9.430 2.800 9.710 3.480 ;
        RECT  11.020 2.800 11.300 3.480 ;
        RECT  11.900 2.800 12.180 3.480 ;
        RECT  13.100 2.800 13.380 3.480 ;
        RECT  14.220 2.800 14.500 3.480 ;
        RECT  15.300 2.620 15.580 3.480 ;
        RECT  16.340 2.620 16.620 3.480 ;
        RECT  17.380 2.620 17.660 3.480 ;
        RECT  18.420 2.620 18.700 3.480 ;
        RECT  0.000 2.920 18.800 3.480 ;
        RECT  0.350 2.800 0.630 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 2.600 8.530 2.760 ;
        RECT  8.370 2.160 8.530 2.760 ;
        RECT  10.930 2.480 15.070 2.640 ;
        RECT  14.910 2.280 15.070 2.640 ;
        RECT  7.180 2.300 7.720 2.640 ;
        RECT  4.420 2.480 7.720 2.640 ;
        RECT  14.440 0.900 14.600 2.640 ;
        RECT  10.930 2.160 11.090 2.640 ;
        RECT  4.420 1.940 4.580 2.640 ;
        RECT  14.910 2.280 16.760 2.440 ;
        RECT  16.600 1.300 16.760 2.440 ;
        RECT  8.370 2.160 11.090 2.320 ;
        RECT  7.560 0.460 7.720 2.760 ;
        RECT  2.540 1.940 4.580 2.100 ;
        RECT  2.540 1.100 2.700 2.100 ;
        RECT  13.980 0.900 14.600 1.060 ;
        RECT  13.980 0.750 14.200 1.060 ;
        RECT  7.400 0.460 7.720 0.680 ;
        RECT  12.460 2.160 14.240 2.320 ;
        RECT  14.080 1.240 14.240 2.320 ;
        RECT  13.660 1.240 14.240 1.400 ;
        RECT  13.660 0.780 13.820 1.400 ;
        RECT  12.560 0.780 12.880 1.040 ;
        RECT  12.560 0.780 13.820 0.940 ;
        RECT  7.880 2.280 8.210 2.440 ;
        RECT  7.880 0.440 8.040 2.440 ;
        RECT  12.780 1.200 12.940 1.940 ;
        RECT  12.200 1.200 12.940 1.360 ;
        RECT  12.200 0.790 12.360 1.360 ;
        RECT  11.360 0.790 12.360 0.950 ;
        RECT  11.360 0.560 11.520 0.950 ;
        RECT  9.670 0.560 11.520 0.720 ;
        RECT  7.880 0.440 9.830 0.600 ;
        RECT  11.250 2.160 11.870 2.320 ;
        RECT  11.250 1.840 11.410 2.320 ;
        RECT  8.780 1.840 11.410 2.000 ;
        RECT  9.780 1.500 11.060 1.660 ;
        RECT  10.900 0.880 11.060 1.660 ;
        RECT  9.780 1.200 9.940 1.660 ;
        RECT  8.720 1.200 9.940 1.360 ;
        RECT  8.720 0.830 8.880 1.360 ;
        RECT  10.900 0.880 11.120 1.160 ;
        RECT  8.780 2.480 10.770 2.640 ;
        RECT  10.160 1.160 10.540 1.320 ;
        RECT  10.160 0.880 10.320 1.320 ;
        RECT  9.140 0.880 10.320 1.040 ;
        RECT  9.140 0.760 9.420 1.040 ;
        RECT  8.200 1.520 8.580 1.980 ;
        RECT  8.200 1.520 9.570 1.680 ;
        RECT  8.200 0.840 8.360 1.980 ;
        RECT  3.980 2.260 4.260 2.520 ;
        RECT  1.660 2.260 4.260 2.420 ;
        RECT  2.220 0.780 2.380 2.420 ;
        RECT  7.240 0.880 7.400 2.040 ;
        RECT  7.080 0.560 7.240 1.040 ;
        RECT  1.590 0.780 3.180 0.940 ;
        RECT  3.020 0.560 3.180 0.940 ;
        RECT  3.020 0.560 7.240 0.720 ;
        RECT  6.760 0.880 6.920 2.320 ;
        RECT  6.760 1.380 7.060 1.660 ;
        RECT  6.700 0.880 6.920 1.160 ;
        RECT  5.540 2.160 6.530 2.320 ;
        RECT  6.370 0.880 6.530 2.320 ;
        RECT  5.540 0.880 6.530 1.040 ;
        RECT  4.920 0.880 5.080 2.320 ;
        RECT  2.910 1.200 3.500 1.360 ;
        RECT  3.340 0.880 3.500 1.360 ;
        RECT  3.340 0.880 5.080 1.040 ;
        RECT  1.320 2.580 2.900 2.740 ;
        RECT  1.320 2.240 1.480 2.740 ;
        RECT  0.820 2.240 1.480 2.400 ;
        RECT  0.860 0.460 1.080 1.020 ;
        RECT  0.860 0.460 2.860 0.620 ;
        RECT  0.440 2.220 0.640 2.500 ;
        RECT  0.480 0.700 0.640 2.500 ;
        RECT  0.480 1.920 2.060 2.080 ;
        RECT  1.900 1.380 2.060 2.080 ;
        RECT  0.380 0.700 0.640 0.980 ;
    END
END DFZERSBKHD

MACRO DFZHHD
    CLASS CORE ;
    FOREIGN DFZHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.350 3.190 1.630 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.960 9.100 2.120 ;
        RECT  8.720 1.840 9.100 2.120 ;
        RECT  8.720 0.960 9.100 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 0.880 10.300 2.120 ;
        RECT  9.840 1.840 10.300 2.120 ;
        RECT  9.840 0.880 10.300 1.160 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 3.330 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  8.100 -0.280 8.380 0.400 ;
        RECT  9.220 -0.280 9.500 0.400 ;
        RECT  10.300 -0.280 10.580 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.520 3.480 ;
        RECT  6.570 2.800 6.850 3.480 ;
        RECT  8.140 2.620 8.420 3.480 ;
        RECT  9.220 2.800 9.500 3.480 ;
        RECT  10.300 2.620 10.580 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  7.700 2.300 11.040 2.460 ;
        RECT  10.880 0.500 11.040 2.460 ;
        RECT  4.240 2.300 4.820 2.460 ;
        RECT  7.300 2.220 7.860 2.380 ;
        RECT  5.490 2.160 6.030 2.320 ;
        RECT  8.400 1.370 8.560 2.460 ;
        RECT  7.300 2.030 7.460 2.380 ;
        RECT  5.870 2.030 7.460 2.190 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  7.620 1.840 8.060 2.060 ;
        RECT  7.900 0.640 8.060 2.060 ;
        RECT  9.520 0.640 9.680 1.710 ;
        RECT  7.780 0.440 7.940 0.970 ;
        RECT  7.780 0.640 9.680 0.800 ;
        RECT  7.500 0.440 7.940 0.600 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.480 1.350 7.700 1.630 ;
        RECT  5.620 1.350 7.700 1.510 ;
        RECT  5.620 0.460 5.780 1.510 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  6.380 0.940 7.460 1.100 ;
        RECT  6.380 0.460 6.540 1.100 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  6.980 2.540 7.460 2.700 ;
        RECT  5.900 2.480 6.430 2.640 ;
        RECT  6.980 2.360 7.140 2.700 ;
        RECT  6.270 2.360 7.140 2.520 ;
        RECT  5.300 1.680 5.700 1.980 ;
        RECT  5.300 1.680 7.280 1.840 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.660 0.560 3.680 0.720 ;
        RECT  3.520 0.440 4.380 0.600 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  3.860 0.760 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.920 3.680 2.310 ;
        RECT  2.760 0.920 3.680 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END DFZHHD

MACRO DFZKHD
    CLASS CORE ;
    FOREIGN DFZKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.780 ;
        RECT  3.260 1.350 3.500 1.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.960 0.960 10.240 1.240 ;
        RECT  9.120 1.840 10.320 2.120 ;
        RECT  9.700 0.960 9.900 2.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.200 0.880 12.400 1.160 ;
        RECT  11.200 1.840 12.400 2.120 ;
        RECT  11.700 0.880 11.900 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.440 -0.280 3.720 0.400 ;
        RECT  6.900 -0.280 7.180 0.420 ;
        RECT  8.340 -0.280 8.620 0.400 ;
        RECT  9.460 -0.280 9.740 0.400 ;
        RECT  10.580 -0.280 10.860 0.400 ;
        RECT  11.660 -0.280 11.940 0.580 ;
        RECT  12.700 -0.280 12.980 0.580 ;
        RECT  0.000 -0.280 13.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.720 3.480 ;
        RECT  7.000 2.800 7.280 3.480 ;
        RECT  8.540 2.620 8.820 3.480 ;
        RECT  9.580 2.620 9.860 3.480 ;
        RECT  10.620 2.620 10.900 3.480 ;
        RECT  11.660 2.620 11.940 3.480 ;
        RECT  12.700 2.620 12.980 3.480 ;
        RECT  0.000 2.920 13.600 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.860 2.600 5.850 2.760 ;
        RECT  5.690 2.160 5.850 2.760 ;
        RECT  4.860 0.460 5.020 2.760 ;
        RECT  8.780 2.300 13.440 2.460 ;
        RECT  13.280 0.500 13.440 2.460 ;
        RECT  4.440 2.300 5.020 2.460 ;
        RECT  7.760 2.280 8.940 2.440 ;
        RECT  5.690 2.160 6.230 2.320 ;
        RECT  8.780 1.400 8.940 2.460 ;
        RECT  7.760 2.000 7.920 2.440 ;
        RECT  6.070 2.000 7.920 2.160 ;
        RECT  4.740 0.460 5.020 0.680 ;
        RECT  8.080 1.840 8.280 2.120 ;
        RECT  8.120 0.640 8.280 2.120 ;
        RECT  10.880 0.640 11.040 1.710 ;
        RECT  7.960 0.640 8.280 0.870 ;
        RECT  7.960 0.640 11.040 0.800 ;
        RECT  7.780 0.440 8.180 0.660 ;
        RECT  5.180 2.180 5.530 2.440 ;
        RECT  5.180 0.460 5.340 2.440 ;
        RECT  7.680 1.260 7.960 1.580 ;
        RECT  5.820 1.260 7.960 1.420 ;
        RECT  5.820 0.460 5.980 1.420 ;
        RECT  5.180 0.460 5.980 0.620 ;
        RECT  7.440 2.600 7.920 2.760 ;
        RECT  6.100 2.480 6.630 2.640 ;
        RECT  7.440 2.340 7.600 2.760 ;
        RECT  6.470 2.340 7.600 2.500 ;
        RECT  6.580 0.940 7.660 1.100 ;
        RECT  6.580 0.460 6.740 1.100 ;
        RECT  6.140 0.460 6.740 0.740 ;
        RECT  5.500 1.580 5.900 1.980 ;
        RECT  5.500 1.580 7.480 1.740 ;
        RECT  5.500 0.840 5.660 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.540 0.880 4.700 2.080 ;
        RECT  4.420 0.560 4.580 1.040 ;
        RECT  1.660 0.560 4.580 0.720 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  4.060 0.880 4.220 2.320 ;
        RECT  4.060 1.380 4.380 1.660 ;
        RECT  4.000 0.880 4.220 1.160 ;
        RECT  2.840 2.150 3.840 2.310 ;
        RECT  3.680 0.920 3.840 2.310 ;
        RECT  3.680 1.460 3.900 1.740 ;
        RECT  2.840 0.920 3.840 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END DFZKHD

MACRO DFZRBCHD
    CLASS CORE ;
    FOREIGN DFZRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 0.840 11.900 2.390 ;
        RECT  11.680 2.110 11.900 2.390 ;
        RECT  11.680 0.840 11.900 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.720 1.240 ;
        RECT  10.500 1.840 10.800 2.120 ;
        RECT  10.500 0.880 10.700 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.540 -0.280 3.820 0.400 ;
        RECT  8.540 -0.280 8.820 0.400 ;
        RECT  9.530 -0.280 9.810 0.400 ;
        RECT  11.060 -0.280 11.340 0.400 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.560 2.800 3.840 3.480 ;
        RECT  8.020 2.800 8.750 3.480 ;
        RECT  9.590 2.800 9.870 3.480 ;
        RECT  11.100 2.280 11.380 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.000 2.600 6.080 2.760 ;
        RECT  5.920 2.140 6.080 2.760 ;
        RECT  7.800 2.480 10.320 2.640 ;
        RECT  10.160 0.440 10.320 2.640 ;
        RECT  5.000 0.460 5.160 2.760 ;
        RECT  7.800 2.140 7.960 2.640 ;
        RECT  4.580 2.300 5.160 2.460 ;
        RECT  5.920 2.140 7.960 2.300 ;
        RECT  11.320 0.560 11.480 1.660 ;
        RECT  10.100 0.560 11.480 0.720 ;
        RECT  4.840 0.460 5.160 0.680 ;
        RECT  10.100 0.440 10.380 0.720 ;
        RECT  8.990 2.160 9.750 2.320 ;
        RECT  9.590 0.980 9.750 2.320 ;
        RECT  9.590 1.460 9.910 1.740 ;
        RECT  5.320 2.220 5.650 2.440 ;
        RECT  5.320 0.440 5.480 2.440 ;
        RECT  9.270 0.620 9.430 1.720 ;
        RECT  8.220 0.620 9.430 0.780 ;
        RECT  8.220 0.440 8.380 0.780 ;
        RECT  5.320 0.440 8.380 0.600 ;
        RECT  8.120 1.820 8.280 2.230 ;
        RECT  6.220 1.820 8.280 1.980 ;
        RECT  7.300 1.080 7.460 1.980 ;
        RECT  7.300 1.080 7.740 1.300 ;
        RECT  6.160 1.080 7.740 1.240 ;
        RECT  6.160 0.840 6.320 1.240 ;
        RECT  7.740 1.460 8.060 1.620 ;
        RECT  7.900 0.760 8.060 1.620 ;
        RECT  6.540 0.760 8.060 0.920 ;
        RECT  7.420 2.460 7.640 2.740 ;
        RECT  6.500 2.460 7.640 2.620 ;
        RECT  5.640 1.400 6.020 1.980 ;
        RECT  5.640 1.400 7.100 1.560 ;
        RECT  5.640 0.840 5.800 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.680 0.880 4.840 2.080 ;
        RECT  4.520 0.520 4.680 1.040 ;
        RECT  1.620 0.560 4.090 0.720 ;
        RECT  3.930 0.520 4.680 0.680 ;
        RECT  4.200 0.840 4.360 2.540 ;
        RECT  4.200 1.380 4.520 1.660 ;
        RECT  2.940 2.320 4.040 2.480 ;
        RECT  3.880 0.880 4.040 2.480 ;
        RECT  2.940 0.880 4.040 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END DFZRBCHD

MACRO DFZRBEHD
    CLASS CORE ;
    FOREIGN DFZRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.280 9.100 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 0.840 11.900 2.390 ;
        RECT  11.680 2.110 11.900 2.390 ;
        RECT  11.680 0.840 11.900 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.000 11.100 2.080 ;
        RECT  10.580 1.880 11.100 2.080 ;
        RECT  10.580 1.000 11.100 1.200 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.710 -0.280 3.990 0.400 ;
        RECT  8.710 -0.280 8.990 0.400 ;
        RECT  9.680 -0.280 9.960 0.400 ;
        RECT  11.100 -0.280 11.380 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.730 2.800 4.010 3.480 ;
        RECT  8.190 2.800 8.920 3.480 ;
        RECT  9.760 2.800 10.040 3.480 ;
        RECT  11.100 2.620 11.380 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.170 2.600 6.250 2.760 ;
        RECT  6.090 2.140 6.250 2.760 ;
        RECT  7.970 2.480 10.460 2.640 ;
        RECT  10.260 2.300 10.460 2.640 ;
        RECT  5.170 0.460 5.330 2.760 ;
        RECT  7.970 2.140 8.130 2.640 ;
        RECT  10.260 2.300 11.480 2.460 ;
        RECT  11.320 1.300 11.480 2.460 ;
        RECT  4.750 2.300 5.330 2.460 ;
        RECT  6.090 2.140 8.130 2.300 ;
        RECT  10.260 0.440 10.420 2.640 ;
        RECT  10.260 0.440 10.460 0.720 ;
        RECT  5.010 0.460 5.330 0.680 ;
        RECT  9.160 2.160 9.920 2.320 ;
        RECT  9.760 0.980 9.920 2.320 ;
        RECT  9.760 1.460 10.080 1.740 ;
        RECT  5.490 2.220 5.820 2.440 ;
        RECT  5.490 0.440 5.650 2.440 ;
        RECT  9.440 0.620 9.600 1.720 ;
        RECT  8.390 0.620 9.600 0.780 ;
        RECT  8.390 0.440 8.550 0.780 ;
        RECT  5.490 0.440 8.550 0.600 ;
        RECT  8.290 1.820 8.450 2.220 ;
        RECT  6.390 1.820 8.450 1.980 ;
        RECT  7.590 1.080 7.750 1.980 ;
        RECT  7.590 1.080 7.910 1.300 ;
        RECT  6.330 1.080 7.910 1.240 ;
        RECT  6.330 0.840 6.490 1.240 ;
        RECT  7.910 1.460 8.230 1.620 ;
        RECT  8.070 0.760 8.230 1.620 ;
        RECT  6.750 0.760 8.230 0.920 ;
        RECT  7.590 2.460 7.810 2.740 ;
        RECT  6.670 2.460 7.810 2.620 ;
        RECT  5.810 1.400 6.190 1.980 ;
        RECT  5.810 1.400 7.280 1.560 ;
        RECT  5.810 0.840 5.970 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.850 0.880 5.010 2.080 ;
        RECT  4.690 0.520 4.850 1.040 ;
        RECT  1.620 0.560 4.260 0.720 ;
        RECT  4.100 0.520 4.850 0.680 ;
        RECT  4.370 0.840 4.530 2.540 ;
        RECT  4.370 1.380 4.690 1.660 ;
        RECT  3.110 2.420 4.210 2.580 ;
        RECT  4.050 0.880 4.210 2.580 ;
        RECT  3.110 0.880 4.210 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.790 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END DFZRBEHD

MACRO DFZRBHHD
    CLASS CORE ;
    FOREIGN DFZRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.440 3.560 1.720 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 0.790 12.700 2.360 ;
        RECT  12.360 2.080 12.700 2.360 ;
        RECT  12.360 0.820 12.700 1.100 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.610 11.500 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.560 -0.280 3.840 0.400 ;
        RECT  8.610 -0.280 8.890 0.400 ;
        RECT  10.740 -0.280 11.020 0.580 ;
        RECT  11.780 -0.280 12.060 0.580 ;
        RECT  12.820 -0.280 13.100 0.580 ;
        RECT  0.000 -0.280 13.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.580 2.800 3.860 3.480 ;
        RECT  8.670 2.740 9.010 3.480 ;
        RECT  9.690 2.620 9.970 3.480 ;
        RECT  10.740 2.620 11.020 3.480 ;
        RECT  11.780 2.620 12.060 3.480 ;
        RECT  12.820 2.620 13.100 3.480 ;
        RECT  0.000 2.920 13.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.020 2.600 8.510 2.760 ;
        RECT  8.350 2.420 8.510 2.760 ;
        RECT  5.020 0.460 5.180 2.760 ;
        RECT  8.350 2.420 9.480 2.580 ;
        RECT  12.040 1.420 12.200 2.460 ;
        RECT  4.600 2.300 5.180 2.460 ;
        RECT  9.320 2.300 12.200 2.460 ;
        RECT  10.240 0.890 10.400 2.460 ;
        RECT  4.860 0.460 5.180 0.680 ;
        RECT  9.130 1.980 9.850 2.140 ;
        RECT  9.690 0.600 9.850 2.140 ;
        RECT  9.690 1.460 10.050 1.740 ;
        RECT  5.340 2.220 5.670 2.440 ;
        RECT  5.340 0.440 5.500 2.440 ;
        RECT  9.370 0.560 9.530 1.680 ;
        RECT  8.220 0.560 9.530 0.720 ;
        RECT  5.340 0.440 8.380 0.600 ;
        RECT  6.610 2.280 8.190 2.440 ;
        RECT  8.030 1.460 8.190 2.440 ;
        RECT  7.640 1.460 8.190 1.620 ;
        RECT  7.900 0.760 8.060 1.620 ;
        RECT  6.560 0.760 8.060 0.920 ;
        RECT  6.920 1.960 7.870 2.120 ;
        RECT  7.590 1.900 7.870 2.120 ;
        RECT  6.240 1.820 7.080 1.980 ;
        RECT  6.920 1.080 7.080 2.120 ;
        RECT  7.460 1.080 7.740 1.300 ;
        RECT  6.180 1.080 7.740 1.240 ;
        RECT  6.180 0.840 6.340 1.240 ;
        RECT  5.660 1.400 6.040 1.980 ;
        RECT  5.660 1.400 6.750 1.560 ;
        RECT  5.660 0.840 5.820 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.700 0.880 4.860 2.040 ;
        RECT  4.540 0.520 4.700 1.040 ;
        RECT  1.610 0.560 4.110 0.720 ;
        RECT  3.950 0.520 4.700 0.680 ;
        RECT  4.220 0.840 4.380 2.540 ;
        RECT  4.220 1.380 4.540 1.660 ;
        RECT  2.960 2.420 4.060 2.580 ;
        RECT  3.900 0.880 4.060 2.580 ;
        RECT  2.960 0.880 4.060 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END DFZRBHHD

MACRO DFZRBKHD
    CLASS CORE ;
    FOREIGN DFZRBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.440 3.560 1.720 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.070 0.860 14.760 1.140 ;
        RECT  13.250 2.060 14.760 2.340 ;
        RECT  13.700 0.860 13.900 2.340 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.970 0.860 12.660 1.140 ;
        RECT  10.970 1.840 12.660 2.120 ;
        RECT  11.700 0.860 11.900 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.560 -0.280 3.840 0.400 ;
        RECT  8.610 -0.280 8.890 0.400 ;
        RECT  10.630 -0.280 10.910 0.580 ;
        RECT  11.690 -0.280 11.970 0.580 ;
        RECT  12.730 -0.280 13.010 0.580 ;
        RECT  13.770 -0.280 14.050 0.580 ;
        RECT  14.810 -0.280 15.090 0.580 ;
        RECT  0.000 -0.280 15.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.580 2.800 3.860 3.480 ;
        RECT  8.670 2.740 10.010 3.480 ;
        RECT  10.630 2.620 10.910 3.480 ;
        RECT  11.690 2.620 11.970 3.480 ;
        RECT  12.730 2.620 13.010 3.480 ;
        RECT  13.770 2.620 14.050 3.480 ;
        RECT  14.810 2.620 15.090 3.480 ;
        RECT  0.000 2.920 15.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.020 2.600 8.510 2.760 ;
        RECT  8.350 2.420 8.510 2.760 ;
        RECT  5.020 0.460 5.180 2.760 ;
        RECT  8.350 2.420 10.370 2.580 ;
        RECT  10.210 0.890 10.370 2.580 ;
        RECT  12.910 1.460 13.070 2.460 ;
        RECT  4.600 2.300 5.180 2.460 ;
        RECT  10.130 2.300 13.070 2.460 ;
        RECT  10.130 1.840 10.370 2.580 ;
        RECT  12.910 1.460 13.130 1.740 ;
        RECT  10.130 0.890 10.370 1.240 ;
        RECT  4.860 0.460 5.180 0.680 ;
        RECT  9.130 2.100 9.850 2.260 ;
        RECT  9.690 0.770 9.850 2.260 ;
        RECT  9.690 1.400 10.050 1.680 ;
        RECT  9.630 0.770 9.850 1.050 ;
        RECT  5.340 2.220 5.670 2.440 ;
        RECT  5.340 0.440 5.500 2.440 ;
        RECT  9.310 1.400 9.530 1.680 ;
        RECT  9.310 0.560 9.470 1.680 ;
        RECT  8.220 0.560 9.470 0.720 ;
        RECT  5.340 0.440 8.380 0.600 ;
        RECT  6.610 2.280 8.190 2.440 ;
        RECT  8.030 1.460 8.190 2.440 ;
        RECT  7.630 1.460 8.190 1.620 ;
        RECT  7.900 0.760 8.060 1.620 ;
        RECT  6.560 0.760 8.060 0.920 ;
        RECT  6.920 1.960 7.870 2.120 ;
        RECT  7.590 1.900 7.870 2.120 ;
        RECT  6.240 1.820 7.080 1.980 ;
        RECT  6.920 1.080 7.080 2.120 ;
        RECT  7.460 1.080 7.740 1.300 ;
        RECT  6.180 1.080 7.740 1.240 ;
        RECT  6.180 0.840 6.340 1.240 ;
        RECT  5.660 1.400 6.040 1.980 ;
        RECT  5.660 1.400 6.740 1.560 ;
        RECT  5.660 0.840 5.820 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.700 0.880 4.860 2.080 ;
        RECT  4.540 0.520 4.700 1.040 ;
        RECT  1.620 0.560 4.110 0.720 ;
        RECT  3.950 0.520 4.700 0.680 ;
        RECT  4.220 0.840 4.380 2.540 ;
        RECT  4.220 1.380 4.540 1.660 ;
        RECT  2.960 2.170 4.060 2.330 ;
        RECT  3.900 0.880 4.060 2.330 ;
        RECT  2.960 0.880 4.060 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END DFZRBKHD

MACRO DFZRSBEHD
    CLASS CORE ;
    FOREIGN DFZRSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.780 0.840 9.100 1.340 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.110 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.420 2.300 1.990 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.080 1.840 12.300 2.120 ;
        RECT  12.100 0.920 12.300 2.160 ;
        RECT  12.080 0.960 12.300 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.960 11.260 1.240 ;
        RECT  10.900 1.840 11.260 2.120 ;
        RECT  10.900 0.960 11.100 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 1.420 9.920 1.700 ;
        RECT  9.700 1.420 9.900 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 -0.280 3.280 0.400 ;
        RECT  7.120 -0.280 7.400 0.620 ;
        RECT  8.560 -0.280 8.840 0.620 ;
        RECT  9.780 -0.280 10.060 0.620 ;
        RECT  11.500 -0.280 11.780 0.580 ;
        RECT  0.000 -0.280 12.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 2.800 2.620 3.480 ;
        RECT  3.160 2.800 3.440 3.480 ;
        RECT  6.620 2.800 6.900 3.480 ;
        RECT  8.220 2.800 8.500 3.480 ;
        RECT  9.380 2.800 9.660 3.480 ;
        RECT  10.400 2.800 10.680 3.480 ;
        RECT  11.500 2.620 11.780 3.480 ;
        RECT  0.000 2.920 12.400 3.480 ;
        RECT  0.560 2.620 0.840 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.580 2.600 5.810 2.760 ;
        RECT  5.650 2.160 5.810 2.760 ;
        RECT  4.580 0.460 4.740 2.760 ;
        RECT  4.200 2.300 4.740 2.460 ;
        RECT  10.580 2.280 11.880 2.440 ;
        RECT  11.720 1.300 11.880 2.440 ;
        RECT  5.650 2.160 10.740 2.320 ;
        RECT  10.580 0.440 10.740 2.440 ;
        RECT  10.580 0.440 10.900 0.750 ;
        RECT  4.420 0.460 4.740 0.680 ;
        RECT  10.240 0.940 10.400 1.460 ;
        RECT  9.440 0.940 10.400 1.100 ;
        RECT  9.910 2.480 10.240 2.740 ;
        RECT  8.740 2.480 10.240 2.640 ;
        RECT  5.210 2.280 5.490 2.440 ;
        RECT  5.250 1.840 5.410 2.440 ;
        RECT  5.250 1.840 6.140 2.000 ;
        RECT  5.980 1.060 6.140 2.000 ;
        RECT  9.180 1.500 9.340 1.920 ;
        RECT  5.980 1.500 9.340 1.660 ;
        RECT  5.560 1.060 6.140 1.220 ;
        RECT  5.560 0.600 5.720 1.220 ;
        RECT  4.940 0.600 5.720 0.760 ;
        RECT  4.940 0.460 5.280 0.760 ;
        RECT  6.300 1.820 9.020 1.980 ;
        RECT  5.970 2.480 8.160 2.640 ;
        RECT  6.410 1.180 7.900 1.340 ;
        RECT  7.740 0.700 7.900 1.340 ;
        RECT  6.410 0.880 6.570 1.340 ;
        RECT  6.300 0.880 6.570 1.160 ;
        RECT  6.730 0.840 7.580 1.000 ;
        RECT  6.730 0.460 6.890 1.000 ;
        RECT  5.910 0.460 6.890 0.620 ;
        RECT  4.900 0.940 5.060 2.080 ;
        RECT  4.900 1.380 5.820 1.660 ;
        RECT  4.900 0.940 5.260 1.100 ;
        RECT  1.360 2.220 1.880 2.380 ;
        RECT  1.720 0.460 1.880 2.380 ;
        RECT  4.260 0.880 4.420 2.040 ;
        RECT  4.100 0.440 4.260 1.040 ;
        RECT  1.720 0.560 3.600 0.720 ;
        RECT  1.640 0.460 1.960 0.620 ;
        RECT  3.440 0.440 4.260 0.600 ;
        RECT  3.780 0.760 3.940 2.340 ;
        RECT  3.780 1.380 4.080 1.660 ;
        RECT  2.680 2.240 3.600 2.400 ;
        RECT  3.440 0.940 3.600 2.400 ;
        RECT  2.680 0.940 3.600 1.100 ;
        RECT  1.020 2.600 1.960 2.760 ;
        RECT  1.020 2.200 1.180 2.760 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END DFZRSBEHD

MACRO DFZRSBHHD
    CLASS CORE ;
    FOREIGN DFZRSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 1.640 9.500 2.140 ;
        RECT  9.280 1.780 9.500 2.060 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.420 3.500 1.960 ;
        RECT  3.260 1.420 3.500 1.700 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.420 2.700 1.990 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.300 0.920 13.500 2.160 ;
        RECT  13.160 1.840 13.500 2.160 ;
        RECT  13.160 0.920 13.500 1.240 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.060 0.960 12.340 1.240 ;
        RECT  12.060 1.840 12.340 2.120 ;
        RECT  12.100 0.960 12.300 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.420 10.700 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.280 2.800 0.400 ;
        RECT  3.310 -0.280 3.590 0.400 ;
        RECT  7.480 -0.280 7.700 0.680 ;
        RECT  9.000 -0.280 9.280 0.620 ;
        RECT  10.320 -0.280 10.600 0.620 ;
        RECT  11.500 -0.280 11.780 0.400 ;
        RECT  12.580 -0.280 12.860 0.580 ;
        RECT  13.620 -0.280 13.900 0.580 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.470 2.800 3.750 3.480 ;
        RECT  6.930 2.800 7.210 3.480 ;
        RECT  8.350 2.800 8.630 3.480 ;
        RECT  9.180 2.800 9.460 3.480 ;
        RECT  10.380 2.800 10.660 3.480 ;
        RECT  11.500 2.800 11.780 3.480 ;
        RECT  12.580 2.620 12.860 3.480 ;
        RECT  13.620 2.620 13.900 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.890 2.600 6.120 2.760 ;
        RECT  5.960 2.160 6.120 2.760 ;
        RECT  8.450 2.480 12.350 2.640 ;
        RECT  12.190 2.280 12.350 2.640 ;
        RECT  4.890 0.460 5.050 2.760 ;
        RECT  11.720 0.900 11.880 2.640 ;
        RECT  8.450 2.160 8.610 2.640 ;
        RECT  4.510 2.300 5.050 2.460 ;
        RECT  12.190 2.280 13.000 2.440 ;
        RECT  12.840 1.300 13.000 2.440 ;
        RECT  5.960 2.160 8.610 2.320 ;
        RECT  11.220 0.900 11.880 1.060 ;
        RECT  11.220 0.750 11.440 1.060 ;
        RECT  4.730 0.460 5.050 0.680 ;
        RECT  9.740 2.160 11.480 2.320 ;
        RECT  11.320 1.240 11.480 2.320 ;
        RECT  10.880 1.240 11.480 1.400 ;
        RECT  10.880 0.780 11.040 1.400 ;
        RECT  9.840 0.780 10.160 1.040 ;
        RECT  9.840 0.780 11.040 0.940 ;
        RECT  5.520 2.280 5.800 2.440 ;
        RECT  5.560 1.840 5.720 2.440 ;
        RECT  5.560 1.840 6.450 2.000 ;
        RECT  6.290 1.060 6.450 2.000 ;
        RECT  10.060 1.200 10.220 1.940 ;
        RECT  6.290 1.500 8.770 1.660 ;
        RECT  8.610 1.200 8.770 1.660 ;
        RECT  8.610 1.200 10.220 1.360 ;
        RECT  5.870 1.060 6.450 1.220 ;
        RECT  5.870 0.600 6.030 1.220 ;
        RECT  5.250 0.600 6.030 0.760 ;
        RECT  5.250 0.460 5.590 0.760 ;
        RECT  8.770 2.100 9.110 2.320 ;
        RECT  8.770 1.820 8.930 2.320 ;
        RECT  6.610 1.820 8.930 1.980 ;
        RECT  7.040 0.840 8.020 1.000 ;
        RECT  7.860 0.560 8.020 1.000 ;
        RECT  7.040 0.460 7.200 1.000 ;
        RECT  7.860 0.560 8.580 0.720 ;
        RECT  6.220 0.460 7.200 0.620 ;
        RECT  6.720 1.180 8.400 1.340 ;
        RECT  8.180 0.880 8.400 1.340 ;
        RECT  6.720 0.880 6.880 1.340 ;
        RECT  6.610 0.880 6.880 1.160 ;
        RECT  6.280 2.480 8.290 2.640 ;
        RECT  5.210 0.940 5.370 2.080 ;
        RECT  5.210 1.380 6.130 1.660 ;
        RECT  5.210 0.940 5.570 1.100 ;
        RECT  1.480 2.520 2.340 2.680 ;
        RECT  2.180 0.560 2.340 2.680 ;
        RECT  4.570 0.880 4.730 2.040 ;
        RECT  4.410 0.440 4.570 1.040 ;
        RECT  1.600 0.740 2.340 0.900 ;
        RECT  2.180 0.560 3.910 0.720 ;
        RECT  3.750 0.440 4.570 0.600 ;
        RECT  4.090 0.760 4.250 2.340 ;
        RECT  4.090 1.380 4.390 1.660 ;
        RECT  2.990 2.180 3.910 2.340 ;
        RECT  3.750 0.880 3.910 2.340 ;
        RECT  2.990 0.880 3.910 1.040 ;
        RECT  0.900 2.200 2.020 2.360 ;
        RECT  1.860 1.460 2.020 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END DFZRSBHHD

MACRO DFZSBEHD
    CLASS CORE ;
    FOREIGN DFZSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.420 3.500 1.960 ;
        RECT  3.270 1.480 3.500 1.760 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.420 2.700 1.990 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.840 11.500 2.260 ;
        RECT  11.280 1.980 11.500 2.260 ;
        RECT  11.280 0.840 11.500 1.120 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.700 2.120 ;
        RECT  10.240 1.840 10.700 2.120 ;
        RECT  10.240 0.960 10.700 1.240 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.260 8.460 1.540 ;
        RECT  8.100 1.140 8.300 1.660 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.280 2.800 0.400 ;
        RECT  3.310 -0.280 3.590 0.400 ;
        RECT  6.990 -0.280 7.270 0.400 ;
        RECT  9.700 -0.280 9.980 0.400 ;
        RECT  10.700 -0.280 10.980 0.580 ;
        RECT  0.000 -0.280 11.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.470 2.800 3.750 3.480 ;
        RECT  6.980 2.800 7.260 3.480 ;
        RECT  7.740 2.800 8.020 3.480 ;
        RECT  8.980 2.800 9.260 3.480 ;
        RECT  10.700 2.620 10.980 3.480 ;
        RECT  0.000 2.920 11.600 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.890 2.600 5.880 2.760 ;
        RECT  5.720 2.160 5.880 2.760 ;
        RECT  6.980 2.480 10.370 2.640 ;
        RECT  10.210 2.300 10.370 2.640 ;
        RECT  4.890 0.460 5.050 2.760 ;
        RECT  8.740 0.940 8.900 2.640 ;
        RECT  6.980 2.160 7.140 2.640 ;
        RECT  10.210 2.300 11.100 2.460 ;
        RECT  10.940 1.460 11.100 2.460 ;
        RECT  4.510 2.300 5.050 2.460 ;
        RECT  5.720 2.160 7.140 2.320 ;
        RECT  10.940 1.460 11.140 1.740 ;
        RECT  8.740 0.940 9.220 1.100 ;
        RECT  4.730 0.460 5.050 0.680 ;
        RECT  9.760 0.650 9.920 2.320 ;
        RECT  9.100 2.150 9.920 2.310 ;
        RECT  9.100 1.620 9.260 2.310 ;
        RECT  9.760 1.400 10.270 1.680 ;
        RECT  5.210 2.280 5.560 2.440 ;
        RECT  5.210 0.460 5.370 2.440 ;
        RECT  9.380 0.440 9.540 1.400 ;
        RECT  5.850 0.900 7.200 1.060 ;
        RECT  7.040 0.560 7.200 1.060 ;
        RECT  5.850 0.460 6.010 1.060 ;
        RECT  7.040 0.560 7.610 0.720 ;
        RECT  5.210 0.460 6.010 0.620 ;
        RECT  7.450 0.440 9.540 0.600 ;
        RECT  7.300 2.060 8.580 2.220 ;
        RECT  8.300 1.920 8.580 2.220 ;
        RECT  7.300 2.000 7.670 2.220 ;
        RECT  7.510 0.880 7.670 2.220 ;
        RECT  6.510 1.360 7.670 1.520 ;
        RECT  7.360 0.880 7.670 1.520 ;
        RECT  5.530 1.680 5.960 1.980 ;
        RECT  5.530 1.680 7.350 1.840 ;
        RECT  5.530 0.840 5.690 1.980 ;
        RECT  6.170 0.460 6.830 0.740 ;
        RECT  6.040 2.480 6.820 2.760 ;
        RECT  1.480 2.520 2.340 2.680 ;
        RECT  2.180 0.560 2.340 2.680 ;
        RECT  4.570 0.880 4.730 2.040 ;
        RECT  4.410 0.440 4.570 1.040 ;
        RECT  1.600 0.740 2.340 0.900 ;
        RECT  2.180 0.560 3.910 0.720 ;
        RECT  3.750 0.440 4.570 0.600 ;
        RECT  4.090 0.760 4.250 2.400 ;
        RECT  4.090 1.380 4.390 1.660 ;
        RECT  3.030 2.240 3.910 2.460 ;
        RECT  3.750 0.880 3.910 2.460 ;
        RECT  3.090 0.880 3.910 1.160 ;
        RECT  0.900 2.200 2.020 2.360 ;
        RECT  1.860 1.460 2.020 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END DFZSBEHD

MACRO DFZSBHHD
    CLASS CORE ;
    FOREIGN DFZSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.420 3.500 1.960 ;
        RECT  3.260 1.480 3.500 1.760 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.420 2.700 1.990 ;
        END
    END TD
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 0.800 12.700 2.360 ;
        RECT  12.360 2.080 12.700 2.360 ;
        RECT  12.360 0.800 12.700 1.080 ;
        END
    END QB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.800 11.500 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.380 8.350 1.660 ;
        RECT  8.100 1.140 8.300 1.660 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.280 2.800 0.400 ;
        RECT  3.300 -0.280 3.580 0.400 ;
        RECT  6.990 -0.280 7.270 0.400 ;
        RECT  8.470 -0.280 8.750 0.400 ;
        RECT  10.700 -0.280 10.980 0.400 ;
        RECT  11.780 -0.280 12.060 0.580 ;
        RECT  12.820 -0.280 13.100 0.580 ;
        RECT  0.000 -0.280 13.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.460 2.800 3.740 3.480 ;
        RECT  7.010 2.800 8.140 3.480 ;
        RECT  8.700 2.800 8.980 3.480 ;
        RECT  9.820 2.800 10.100 3.480 ;
        RECT  10.740 2.620 11.020 3.480 ;
        RECT  11.780 2.620 12.060 3.480 ;
        RECT  12.820 2.620 13.100 3.480 ;
        RECT  0.000 2.920 13.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.880 2.600 5.870 2.760 ;
        RECT  5.710 2.160 5.870 2.760 ;
        RECT  6.990 2.480 9.480 2.640 ;
        RECT  9.320 1.020 9.480 2.640 ;
        RECT  4.880 0.460 5.040 2.760 ;
        RECT  6.990 2.160 7.150 2.640 ;
        RECT  4.500 2.300 5.040 2.460 ;
        RECT  9.320 2.280 12.200 2.440 ;
        RECT  12.040 1.400 12.200 2.440 ;
        RECT  5.710 2.160 7.150 2.320 ;
        RECT  9.320 1.020 9.740 1.180 ;
        RECT  4.720 0.460 5.040 0.680 ;
        RECT  10.180 1.960 11.140 2.120 ;
        RECT  10.980 1.400 11.140 2.120 ;
        RECT  10.180 0.960 10.340 2.120 ;
        RECT  10.020 0.960 10.340 1.620 ;
        RECT  5.200 2.280 5.550 2.440 ;
        RECT  5.200 0.460 5.360 2.440 ;
        RECT  10.500 0.640 10.660 1.620 ;
        RECT  5.840 0.900 7.170 1.060 ;
        RECT  7.010 0.560 7.170 1.060 ;
        RECT  5.840 0.460 6.000 1.060 ;
        RECT  10.200 0.640 10.660 0.800 ;
        RECT  7.010 0.560 10.360 0.720 ;
        RECT  5.200 0.460 6.000 0.620 ;
        RECT  7.310 1.980 7.680 2.280 ;
        RECT  7.520 0.940 7.680 2.280 ;
        RECT  7.310 1.980 8.630 2.140 ;
        RECT  6.520 1.220 6.840 1.480 ;
        RECT  6.520 1.220 7.750 1.380 ;
        RECT  7.470 0.940 7.750 1.380 ;
        RECT  5.520 1.660 5.950 1.980 ;
        RECT  5.520 1.660 7.360 1.820 ;
        RECT  7.080 1.540 7.360 1.820 ;
        RECT  5.520 0.840 5.680 1.980 ;
        RECT  6.250 2.480 6.790 2.760 ;
        RECT  6.180 0.460 6.780 0.740 ;
        RECT  1.480 2.520 2.340 2.680 ;
        RECT  2.180 0.560 2.340 2.680 ;
        RECT  4.560 0.880 4.720 2.040 ;
        RECT  4.400 0.440 4.560 1.040 ;
        RECT  1.600 0.740 2.340 0.900 ;
        RECT  2.180 0.560 3.900 0.720 ;
        RECT  3.740 0.440 4.560 0.600 ;
        RECT  4.080 0.760 4.240 2.450 ;
        RECT  4.080 1.380 4.380 1.660 ;
        RECT  2.980 2.180 3.900 2.340 ;
        RECT  3.740 0.910 3.900 2.340 ;
        RECT  2.980 0.910 3.900 1.070 ;
        RECT  0.900 2.200 2.020 2.360 ;
        RECT  1.860 1.460 2.020 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END DFZSBHHD

MACRO DFZTRBCHD
    CLASS CORE ;
    FOREIGN DFZTRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 0.870 11.900 2.250 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        RECT  8.480 1.400 8.700 1.680 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.410 3.260 1.690 ;
        RECT  2.900 1.240 3.100 1.910 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        END
    END TD
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.500 0.840 12.700 1.560 ;
        RECT  12.480 1.140 12.700 1.420 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.700 2.120 ;
        RECT  10.300 1.840 10.700 2.120 ;
        RECT  10.300 0.960 10.700 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 1.980 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.330 -0.280 3.610 0.400 ;
        RECT  8.290 -0.280 8.570 0.400 ;
        RECT  9.280 -0.280 9.560 0.400 ;
        RECT  10.800 -0.280 11.080 0.580 ;
        RECT  12.120 -0.280 12.400 0.400 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.480 2.800 2.760 3.480 ;
        RECT  3.330 2.800 3.610 3.480 ;
        RECT  7.770 2.800 8.500 3.480 ;
        RECT  9.340 2.800 9.620 3.480 ;
        RECT  10.800 2.620 11.080 3.480 ;
        RECT  12.150 2.800 12.430 3.480 ;
        RECT  0.000 2.920 12.800 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  12.120 1.620 12.340 2.280 ;
        RECT  12.120 0.700 12.280 2.280 ;
        RECT  12.120 0.700 12.340 0.980 ;
        RECT  4.750 2.600 5.830 2.760 ;
        RECT  5.670 2.140 5.830 2.760 ;
        RECT  7.550 2.480 10.120 2.640 ;
        RECT  9.850 2.350 10.120 2.640 ;
        RECT  4.750 0.460 4.910 2.760 ;
        RECT  7.550 2.140 7.710 2.640 ;
        RECT  4.330 2.300 4.910 2.460 ;
        RECT  9.850 0.460 10.010 2.640 ;
        RECT  5.670 2.140 7.710 2.300 ;
        RECT  9.850 0.460 10.070 0.740 ;
        RECT  4.590 0.460 4.910 0.680 ;
        RECT  8.740 2.160 9.500 2.320 ;
        RECT  9.340 0.980 9.500 2.320 ;
        RECT  9.340 1.460 9.660 1.740 ;
        RECT  5.070 2.220 5.400 2.440 ;
        RECT  5.070 0.440 5.230 2.440 ;
        RECT  9.020 0.620 9.180 1.720 ;
        RECT  7.970 0.620 9.180 0.780 ;
        RECT  7.970 0.440 8.130 0.780 ;
        RECT  5.070 0.440 8.130 0.600 ;
        RECT  7.870 1.820 8.030 2.230 ;
        RECT  5.970 1.820 8.030 1.980 ;
        RECT  7.050 1.080 7.210 1.980 ;
        RECT  7.050 1.080 7.490 1.300 ;
        RECT  5.910 1.080 7.490 1.240 ;
        RECT  5.910 0.840 6.070 1.240 ;
        RECT  7.490 1.460 7.810 1.620 ;
        RECT  7.650 0.760 7.810 1.620 ;
        RECT  6.290 0.760 7.810 0.920 ;
        RECT  7.170 2.460 7.390 2.740 ;
        RECT  6.250 2.460 7.390 2.620 ;
        RECT  5.390 1.400 5.770 1.980 ;
        RECT  5.390 1.400 6.850 1.560 ;
        RECT  5.390 0.840 5.550 1.980 ;
        RECT  1.520 2.280 1.880 2.440 ;
        RECT  1.720 0.560 1.880 2.440 ;
        RECT  4.430 0.880 4.590 2.080 ;
        RECT  4.270 0.560 4.430 1.040 ;
        RECT  1.620 0.560 4.430 0.720 ;
        RECT  3.950 0.880 4.110 2.440 ;
        RECT  3.950 1.380 4.270 1.660 ;
        RECT  3.890 0.880 4.110 1.160 ;
        RECT  2.850 2.130 3.730 2.290 ;
        RECT  3.570 0.880 3.730 2.290 ;
        RECT  3.570 1.440 3.790 1.720 ;
        RECT  2.850 0.880 3.730 1.040 ;
        RECT  1.110 2.600 2.200 2.760 ;
        RECT  2.040 1.760 2.200 2.760 ;
        RECT  1.110 2.300 1.270 2.760 ;
        RECT  0.100 2.300 1.270 2.460 ;
        RECT  0.920 1.090 1.080 2.460 ;
        RECT  0.100 2.000 0.320 2.460 ;
        RECT  2.040 1.760 2.260 2.040 ;
        RECT  0.100 0.460 0.260 2.460 ;
        RECT  0.100 0.460 0.380 0.680 ;
    END
END DFZTRBCHD

MACRO DFZTRBEHD
    CLASS CORE ;
    FOREIGN DFZTRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QZ
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.900 0.840 13.100 2.360 ;
        RECT  12.740 2.060 13.100 2.360 ;
        RECT  12.740 0.840 13.100 1.140 ;
        END
    END QZ
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        RECT  8.480 1.400 8.700 1.680 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.410 3.260 1.690 ;
        RECT  2.900 1.240 3.100 1.910 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        END
    END TD
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.100 1.140 14.300 1.860 ;
        RECT  14.080 1.140 14.300 1.420 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.700 2.120 ;
        RECT  10.380 1.840 10.700 2.120 ;
        RECT  10.380 0.960 10.700 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 1.980 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.330 -0.280 3.610 0.400 ;
        RECT  8.290 -0.280 8.570 0.400 ;
        RECT  9.340 -0.280 9.620 0.400 ;
        RECT  10.840 -0.280 11.120 0.580 ;
        RECT  11.880 -0.280 12.160 0.580 ;
        RECT  13.800 -0.280 14.080 0.400 ;
        RECT  0.000 -0.280 14.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.480 2.800 2.760 3.480 ;
        RECT  3.330 2.800 3.610 3.480 ;
        RECT  7.770 2.800 8.500 3.480 ;
        RECT  9.340 2.800 9.620 3.480 ;
        RECT  10.840 2.620 11.120 3.480 ;
        RECT  11.880 2.620 12.160 3.480 ;
        RECT  13.770 2.800 14.050 3.480 ;
        RECT  0.000 2.920 14.400 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  13.720 2.000 13.960 2.280 ;
        RECT  13.720 0.800 13.880 2.280 ;
        RECT  13.720 0.800 14.020 0.960 ;
        RECT  13.320 0.520 13.480 1.130 ;
        RECT  11.310 0.920 12.500 1.080 ;
        RECT  12.340 0.520 12.500 1.080 ;
        RECT  12.340 0.520 13.480 0.680 ;
        RECT  12.340 2.520 13.480 2.680 ;
        RECT  13.320 2.050 13.480 2.680 ;
        RECT  12.340 2.120 12.500 2.680 ;
        RECT  11.310 2.120 12.500 2.280 ;
        RECT  4.750 2.600 5.830 2.760 ;
        RECT  5.670 2.140 5.830 2.760 ;
        RECT  7.550 2.480 10.120 2.640 ;
        RECT  9.960 0.520 10.120 2.640 ;
        RECT  4.750 0.460 4.910 2.760 ;
        RECT  7.550 2.140 7.710 2.640 ;
        RECT  4.330 2.300 4.910 2.460 ;
        RECT  5.670 2.140 7.710 2.300 ;
        RECT  9.900 0.520 10.120 0.800 ;
        RECT  4.590 0.460 4.910 0.680 ;
        RECT  8.740 2.160 9.500 2.320 ;
        RECT  9.340 0.980 9.500 2.320 ;
        RECT  9.340 1.460 9.660 1.740 ;
        RECT  5.070 2.220 5.400 2.440 ;
        RECT  5.070 0.440 5.230 2.440 ;
        RECT  9.020 0.620 9.180 1.720 ;
        RECT  7.970 0.620 9.180 0.780 ;
        RECT  7.970 0.440 8.130 0.780 ;
        RECT  5.070 0.440 8.130 0.600 ;
        RECT  7.870 1.820 8.030 2.230 ;
        RECT  5.970 1.820 8.030 1.980 ;
        RECT  7.050 1.080 7.210 1.980 ;
        RECT  7.050 1.080 7.490 1.300 ;
        RECT  5.910 1.080 7.490 1.240 ;
        RECT  5.910 0.840 6.070 1.240 ;
        RECT  7.490 1.460 7.810 1.620 ;
        RECT  7.650 0.760 7.810 1.620 ;
        RECT  6.290 0.760 7.810 0.920 ;
        RECT  7.170 2.460 7.390 2.740 ;
        RECT  6.250 2.460 7.390 2.620 ;
        RECT  5.390 1.400 5.770 1.980 ;
        RECT  5.390 1.400 6.850 1.560 ;
        RECT  5.390 0.840 5.550 1.980 ;
        RECT  1.520 2.280 1.880 2.440 ;
        RECT  1.720 0.560 1.880 2.440 ;
        RECT  4.430 0.880 4.590 2.080 ;
        RECT  4.270 0.560 4.430 1.040 ;
        RECT  1.620 0.560 4.430 0.720 ;
        RECT  3.950 0.880 4.110 2.440 ;
        RECT  3.950 1.380 4.270 1.660 ;
        RECT  3.890 0.880 4.110 1.160 ;
        RECT  2.850 2.130 3.730 2.290 ;
        RECT  3.570 0.880 3.730 2.290 ;
        RECT  3.570 1.440 3.790 1.720 ;
        RECT  2.850 0.880 3.730 1.040 ;
        RECT  1.110 2.600 2.200 2.760 ;
        RECT  2.040 1.760 2.200 2.760 ;
        RECT  1.110 2.300 1.270 2.760 ;
        RECT  0.100 2.300 1.270 2.460 ;
        RECT  0.920 1.090 1.080 2.460 ;
        RECT  0.100 2.000 0.320 2.460 ;
        RECT  2.040 1.760 2.260 2.040 ;
        RECT  0.100 0.460 0.260 2.460 ;
        RECT  0.100 0.460 0.380 0.680 ;
    END
END DFZTRBEHD

MACRO DLAHCHD
    CLASS CORE ;
    FOREIGN DLAHCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.720 6.700 2.400 ;
        RECT  6.470 2.120 6.700 2.400 ;
        RECT  6.470 0.720 6.700 1.000 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.850 5.510 1.130 ;
        RECT  5.300 1.840 5.510 2.120 ;
        RECT  5.300 0.850 5.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.600 ;
        RECT  5.890 -0.280 6.170 0.940 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.850 2.800 6.130 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 2.300 6.210 2.460 ;
        RECT  6.050 1.420 6.210 2.460 ;
        RECT  4.870 0.440 5.030 2.460 ;
        RECT  4.090 0.860 4.250 1.140 ;
        RECT  4.090 0.920 5.030 1.080 ;
        RECT  4.810 0.440 5.090 0.600 ;
        RECT  3.050 2.480 4.630 2.640 ;
        RECT  4.470 1.460 4.630 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.440 3.850 2.320 ;
        RECT  3.690 0.440 3.970 0.600 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  1.290 0.580 2.370 0.740 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  0.100 2.300 2.870 2.460 ;
        RECT  2.710 1.380 2.870 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.330 1.840 2.550 2.120 ;
        RECT  2.390 0.940 2.550 2.120 ;
        RECT  2.330 0.940 2.610 1.100 ;
    END
END DLAHCHD

MACRO DLAHEHD
    CLASS CORE ;
    FOREIGN DLAHEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.520 6.700 2.680 ;
        RECT  6.470 2.400 6.700 2.680 ;
        RECT  6.470 0.720 6.700 1.000 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.850 5.510 1.130 ;
        RECT  5.300 1.840 5.510 2.120 ;
        RECT  5.300 0.850 5.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.980 ;
        RECT  5.890 -0.280 6.170 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.850 2.800 6.130 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 2.300 6.210 2.460 ;
        RECT  6.050 1.420 6.210 2.460 ;
        RECT  4.870 0.820 5.030 2.460 ;
        RECT  4.030 1.200 4.310 1.420 ;
        RECT  4.030 1.200 5.090 1.360 ;
        RECT  4.810 0.820 5.090 1.360 ;
        RECT  3.050 2.480 4.630 2.640 ;
        RECT  4.470 1.690 4.630 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.820 3.850 2.320 ;
        RECT  3.690 0.820 3.970 0.980 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  1.290 0.580 2.370 0.740 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  0.100 2.300 2.870 2.460 ;
        RECT  2.710 1.380 2.870 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.390 0.940 2.550 2.130 ;
        RECT  2.330 1.850 2.550 2.120 ;
        RECT  2.330 0.940 2.610 1.100 ;
    END
END DLAHEHD

MACRO DLAHHHD
    CLASS CORE ;
    FOREIGN DLAHHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.720 7.150 1.000 ;
        RECT  6.900 2.400 7.150 2.680 ;
        RECT  6.900 0.520 7.100 2.680 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.850 6.030 1.130 ;
        RECT  5.700 1.840 6.030 2.120 ;
        RECT  5.700 0.850 5.900 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.980 ;
        RECT  5.290 -0.280 5.570 0.580 ;
        RECT  6.410 -0.280 6.690 0.580 ;
        RECT  7.530 -0.280 7.810 0.580 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.290 2.620 5.570 3.480 ;
        RECT  6.370 2.620 6.650 3.480 ;
        RECT  7.490 2.620 7.770 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 2.300 6.730 2.460 ;
        RECT  6.570 1.380 6.730 2.460 ;
        RECT  4.870 0.820 5.030 2.460 ;
        RECT  4.030 1.200 4.310 1.420 ;
        RECT  4.030 1.200 5.090 1.360 ;
        RECT  4.810 0.820 5.090 1.360 ;
        RECT  3.050 2.480 4.700 2.640 ;
        RECT  4.540 1.520 4.700 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.820 3.850 2.320 ;
        RECT  3.690 0.820 3.970 0.980 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  1.290 0.580 2.370 0.740 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  0.100 2.300 2.890 2.460 ;
        RECT  2.730 1.440 2.890 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 2.220 0.380 2.460 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.330 1.840 2.550 2.120 ;
        RECT  2.390 0.960 2.550 2.120 ;
    END
END DLAHHHD

MACRO DLAHRBCHD
    CLASS CORE ;
    FOREIGN DLAHRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.340 2.300 1.620 ;
        RECT  2.100 1.000 2.300 1.620 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.720 7.500 2.400 ;
        RECT  7.270 2.120 7.500 2.400 ;
        RECT  7.270 0.720 7.500 1.000 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.340 2.840 1.620 ;
        RECT  2.500 1.000 2.700 1.620 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.850 6.310 1.130 ;
        RECT  6.100 1.840 6.310 2.120 ;
        RECT  6.100 0.850 6.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.660 ;
        RECT  6.690 -0.280 6.970 0.940 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.490 2.470 2.770 3.480 ;
        RECT  5.220 2.740 5.870 3.480 ;
        RECT  6.650 2.800 6.930 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.670 2.300 7.010 2.460 ;
        RECT  6.850 1.420 7.010 2.460 ;
        RECT  5.670 0.440 5.830 2.460 ;
        RECT  4.890 0.940 5.110 1.220 ;
        RECT  4.890 1.000 5.830 1.160 ;
        RECT  2.930 2.600 5.060 2.760 ;
        RECT  4.900 2.420 5.060 2.760 ;
        RECT  3.890 0.820 4.050 2.760 ;
        RECT  2.930 2.150 3.090 2.760 ;
        RECT  4.900 2.420 5.430 2.580 ;
        RECT  5.270 1.460 5.430 2.580 ;
        RECT  1.930 2.150 2.210 2.370 ;
        RECT  1.930 2.150 3.090 2.310 ;
        RECT  3.710 0.820 4.050 0.980 ;
        RECT  4.530 2.130 4.740 2.440 ;
        RECT  4.530 0.440 4.690 2.440 ;
        RECT  4.530 0.440 4.750 0.720 ;
        RECT  1.290 0.560 1.450 2.120 ;
        RECT  4.210 0.440 4.370 2.060 ;
        RECT  1.290 0.560 2.490 0.720 ;
        RECT  2.330 0.440 4.370 0.600 ;
        RECT  3.270 2.150 3.730 2.310 ;
        RECT  3.570 1.140 3.730 2.310 ;
        RECT  3.350 1.140 3.730 1.300 ;
        RECT  3.350 0.820 3.510 1.300 ;
        RECT  3.230 0.820 3.510 1.040 ;
        RECT  0.100 2.300 1.770 2.460 ;
        RECT  1.610 1.830 1.770 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  1.610 1.830 3.410 1.990 ;
        RECT  3.250 1.510 3.410 1.990 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END DLAHRBCHD

MACRO DLAHRBEHD
    CLASS CORE ;
    FOREIGN DLAHRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.340 2.300 1.620 ;
        RECT  2.100 1.000 2.300 1.620 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.520 7.500 2.670 ;
        RECT  7.270 2.390 7.500 2.670 ;
        RECT  7.270 0.520 7.500 0.800 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.340 2.840 1.620 ;
        RECT  2.500 1.000 2.700 1.620 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.850 6.310 1.130 ;
        RECT  6.100 1.840 6.310 2.120 ;
        RECT  6.100 0.850 6.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.760 ;
        RECT  6.690 -0.280 6.970 0.580 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.490 2.470 2.770 3.480 ;
        RECT  5.220 2.740 5.420 3.480 ;
        RECT  6.650 2.800 6.930 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.670 2.300 7.010 2.460 ;
        RECT  6.850 1.420 7.010 2.460 ;
        RECT  5.670 0.540 5.830 2.460 ;
        RECT  4.890 1.070 5.050 1.350 ;
        RECT  4.890 1.130 5.830 1.290 ;
        RECT  2.930 2.600 5.060 2.760 ;
        RECT  4.900 2.420 5.060 2.760 ;
        RECT  3.890 0.820 4.050 2.760 ;
        RECT  2.930 2.150 3.090 2.760 ;
        RECT  4.900 2.420 5.430 2.580 ;
        RECT  5.270 1.550 5.430 2.580 ;
        RECT  1.930 2.150 2.210 2.370 ;
        RECT  1.930 2.150 3.090 2.310 ;
        RECT  3.710 0.820 4.050 0.980 ;
        RECT  4.530 2.130 4.740 2.440 ;
        RECT  4.530 0.540 4.690 2.440 ;
        RECT  1.290 0.560 1.450 2.120 ;
        RECT  4.210 0.440 4.370 2.060 ;
        RECT  1.290 0.560 2.490 0.720 ;
        RECT  2.330 0.440 4.370 0.600 ;
        RECT  3.270 2.150 3.730 2.310 ;
        RECT  3.570 1.140 3.730 2.310 ;
        RECT  3.350 1.140 3.730 1.300 ;
        RECT  3.350 0.820 3.510 1.300 ;
        RECT  3.230 0.820 3.510 1.040 ;
        RECT  0.100 2.300 1.770 2.460 ;
        RECT  1.610 1.830 1.770 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  1.610 1.830 3.410 1.990 ;
        RECT  3.250 1.510 3.410 1.990 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END DLAHRBEHD

MACRO DLAHRBHHD
    CLASS CORE ;
    FOREIGN DLAHRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.000 2.300 1.650 ;
        END
    END RB
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 0.900 8.300 2.300 ;
        RECT  7.820 2.100 8.300 2.300 ;
        RECT  7.820 0.900 8.300 1.100 ;
        END
    END QB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.370 2.970 1.650 ;
        RECT  2.500 1.000 2.700 1.650 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.850 7.100 2.120 ;
        RECT  6.760 1.840 7.100 2.120 ;
        RECT  6.760 0.850 7.100 1.130 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.980 ;
        RECT  6.180 -0.280 6.460 0.580 ;
        RECT  7.300 -0.280 7.580 0.580 ;
        RECT  8.420 -0.280 8.700 0.580 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.620 2.800 3.480 ;
        RECT  5.240 2.320 5.460 3.480 ;
        RECT  6.180 2.620 6.460 3.480 ;
        RECT  7.260 2.620 7.540 3.480 ;
        RECT  8.380 2.620 8.660 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.760 2.300 7.620 2.460 ;
        RECT  7.460 1.420 7.620 2.460 ;
        RECT  5.760 0.820 5.920 2.460 ;
        RECT  4.890 1.140 5.110 1.420 ;
        RECT  4.890 1.200 5.920 1.360 ;
        RECT  5.700 0.820 5.980 0.980 ;
        RECT  2.970 2.600 5.080 2.760 ;
        RECT  4.920 1.940 5.080 2.760 ;
        RECT  3.930 0.760 4.090 2.760 ;
        RECT  2.970 2.300 3.130 2.760 ;
        RECT  1.930 2.300 3.130 2.460 ;
        RECT  4.920 1.940 5.590 2.100 ;
        RECT  5.430 1.520 5.590 2.100 ;
        RECT  4.570 2.130 4.760 2.440 ;
        RECT  4.570 0.760 4.730 2.440 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  4.250 0.440 4.410 2.070 ;
        RECT  1.290 0.580 2.490 0.740 ;
        RECT  2.330 0.440 4.410 0.600 ;
        RECT  3.310 2.240 3.770 2.400 ;
        RECT  3.610 0.940 3.770 2.400 ;
        RECT  3.190 0.940 3.770 1.100 ;
        RECT  3.190 0.820 3.470 1.100 ;
        RECT  0.100 2.300 1.770 2.460 ;
        RECT  1.610 1.920 1.770 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 2.220 0.380 2.460 ;
        RECT  1.610 1.920 3.450 2.080 ;
        RECT  3.290 1.480 3.450 2.080 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END DLAHRBHHD

MACRO FA1DHD
    CLASS CORE ;
    FOREIGN FA1DHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.400 1.080 3.560 1.680 ;
        RECT  3.400 1.520 3.900 1.680 ;
        RECT  3.700 1.520 3.900 2.120 ;
        RECT  3.700 1.960 4.060 2.120 ;
        RECT  3.280 1.080 3.560 1.240 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.600 1.720 1.760 2.760 ;
        RECT  2.410 2.260 2.570 2.760 ;
        RECT  1.600 2.600 2.570 2.760 ;
        RECT  2.410 2.260 3.380 2.420 ;
        RECT  3.220 2.260 3.380 2.600 ;
        RECT  4.520 1.960 4.680 2.600 ;
        RECT  3.220 2.440 4.680 2.600 ;
        RECT  6.740 1.520 7.100 1.800 ;
        RECT  6.900 1.520 7.100 2.120 ;
        RECT  4.520 1.960 7.100 2.120 ;
        RECT  1.460 1.720 1.760 1.940 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.520 8.700 2.280 ;
        RECT  8.480 2.000 8.700 2.280 ;
        RECT  8.480 0.520 8.700 0.800 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 0.620 2.370 0.780 ;
        RECT  2.210 0.760 3.880 0.920 ;
        RECT  3.720 0.760 3.880 1.360 ;
        RECT  3.720 1.200 7.500 1.360 ;
        RECT  7.300 1.200 7.500 1.840 ;
        RECT  1.760 0.440 2.040 0.780 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.340 1.020 1.620 ;
        RECT  0.500 1.240 0.700 1.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 -0.280 2.360 0.460 ;
        RECT  4.360 -0.280 4.520 0.670 ;
        RECT  5.420 -0.280 5.700 0.400 ;
        RECT  7.860 -0.280 8.140 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.160 -0.280 0.320 1.000 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.780 2.580 3.060 3.480 ;
        RECT  4.260 2.790 4.540 3.480 ;
        RECT  5.420 2.800 5.700 3.480 ;
        RECT  7.860 2.800 8.140 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.500 2.300 8.320 2.460 ;
        RECT  8.160 0.560 8.320 2.460 ;
        RECT  8.120 1.340 8.340 1.620 ;
        RECT  6.500 0.560 8.320 0.720 ;
        RECT  7.700 0.880 7.860 1.620 ;
        RECT  4.040 0.880 7.860 1.040 ;
        RECT  4.040 0.440 4.200 1.040 ;
        RECT  2.640 0.440 4.200 0.600 ;
        RECT  6.180 1.520 6.340 1.800 ;
        RECT  4.090 1.520 6.340 1.680 ;
        RECT  4.860 0.560 6.260 0.720 ;
        RECT  4.860 2.480 6.260 2.640 ;
        RECT  5.980 2.280 6.260 2.640 ;
        RECT  1.920 1.400 2.080 2.380 ;
        RECT  1.920 1.520 3.120 1.680 ;
        RECT  1.260 1.400 2.080 1.560 ;
        RECT  1.260 0.740 1.420 1.560 ;
        RECT  1.020 0.740 1.420 0.900 ;
        RECT  1.580 1.080 3.020 1.240 ;
        RECT  1.580 1.020 1.860 1.240 ;
        RECT  1.280 2.420 1.440 2.700 ;
        RECT  0.100 2.480 1.440 2.640 ;
    END
END FA1DHD

MACRO FA1EHD
    CLASS CORE ;
    FOREIGN FA1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  12.480 0.520 12.700 2.280 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.100 0.560 4.780 0.720 ;
        RECT  4.620 0.560 4.780 2.280 ;
        RECT  4.620 2.120 5.100 2.280 ;
        RECT  4.940 2.120 5.100 2.760 ;
        RECT  4.940 2.600 8.180 2.760 ;
        RECT  8.020 2.480 9.070 2.640 ;
        RECT  8.910 2.100 9.070 2.640 ;
        RECT  10.450 1.840 10.610 2.260 ;
        RECT  8.910 2.100 10.610 2.260 ;
        RECT  11.250 1.340 11.500 2.000 ;
        RECT  10.450 1.840 11.500 2.000 ;
        RECT  2.100 0.440 3.260 0.600 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 0.680 0.320 0.960 ;
        RECT  0.100 2.230 0.320 2.510 ;
        RECT  0.100 0.680 0.300 2.510 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.640 1.460 7.920 1.680 ;
        RECT  7.640 1.520 10.320 1.680 ;
        RECT  7.700 1.140 7.900 1.680 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 1.140 10.700 1.660 ;
        RECT  10.500 1.400 10.960 1.560 ;
        RECT  8.320 1.200 10.700 1.360 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.520 -0.280 3.800 0.400 ;
        RECT  5.020 -0.280 5.300 0.400 ;
        RECT  7.880 -0.280 8.040 0.460 ;
        RECT  8.920 -0.280 9.080 0.700 ;
        RECT  9.940 -0.280 10.220 0.400 ;
        RECT  11.860 -0.280 12.140 0.400 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.520 2.800 3.800 3.480 ;
        RECT  4.620 2.740 4.780 3.480 ;
        RECT  8.380 2.800 9.100 3.480 ;
        RECT  9.940 2.800 10.220 3.480 ;
        RECT  11.860 2.800 12.140 3.480 ;
        RECT  0.000 2.920 12.800 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.820 2.160 12.300 2.320 ;
        RECT  12.140 0.880 12.300 2.320 ;
        RECT  10.860 0.880 12.300 1.040 ;
        RECT  9.380 0.560 11.660 0.720 ;
        RECT  9.380 2.480 11.660 2.640 ;
        RECT  5.260 2.280 7.860 2.440 ;
        RECT  7.700 2.000 7.860 2.440 ;
        RECT  6.740 1.960 7.060 2.440 ;
        RECT  5.260 1.250 5.420 2.440 ;
        RECT  7.700 2.000 8.660 2.160 ;
        RECT  6.740 0.440 6.900 2.440 ;
        RECT  5.260 1.250 5.580 1.530 ;
        RECT  7.560 0.730 8.660 0.890 ;
        RECT  7.560 0.440 7.720 0.890 ;
        RECT  6.740 0.440 7.720 0.600 ;
        RECT  7.240 1.840 7.540 2.060 ;
        RECT  7.240 0.760 7.400 2.060 ;
        RECT  7.180 1.320 7.400 1.600 ;
        RECT  6.180 1.960 6.460 2.120 ;
        RECT  6.300 0.560 6.460 2.120 ;
        RECT  4.940 0.560 5.100 1.650 ;
        RECT  6.100 0.880 6.460 1.100 ;
        RECT  4.940 0.560 6.460 0.720 ;
        RECT  5.580 1.840 5.900 2.060 ;
        RECT  5.740 0.880 5.900 2.060 ;
        RECT  5.540 0.880 5.900 1.040 ;
        RECT  1.980 2.480 4.300 2.640 ;
        RECT  4.140 0.880 4.300 2.640 ;
        RECT  1.980 1.080 2.140 2.640 ;
        RECT  3.340 1.380 4.300 1.540 ;
        RECT  1.770 1.080 2.140 1.300 ;
        RECT  1.760 1.080 2.140 1.240 ;
        RECT  3.020 0.880 3.180 2.320 ;
        RECT  2.500 0.760 2.660 2.320 ;
        RECT  0.500 0.560 0.660 1.660 ;
        RECT  1.760 0.760 2.660 0.920 ;
        RECT  1.760 0.560 1.920 0.920 ;
        RECT  0.500 0.560 1.920 0.720 ;
        RECT  1.280 2.020 1.580 2.300 ;
        RECT  1.420 1.020 1.580 2.300 ;
        RECT  1.220 1.020 1.580 1.180 ;
    END
END FA1EHD

MACRO FA1HHD
    CLASS CORE ;
    FOREIGN FA1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.700 0.900 13.900 2.300 ;
        RECT  13.100 2.100 13.900 2.300 ;
        RECT  13.100 0.900 13.900 1.100 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.790 0.560 5.420 0.720 ;
        RECT  5.260 0.560 5.420 2.280 ;
        RECT  5.260 2.120 5.740 2.280 ;
        RECT  5.580 2.120 5.740 2.760 ;
        RECT  8.660 2.360 8.820 2.760 ;
        RECT  5.580 2.600 8.820 2.760 ;
        RECT  9.590 2.100 9.750 2.520 ;
        RECT  8.660 2.360 9.750 2.520 ;
        RECT  11.180 1.840 11.340 2.260 ;
        RECT  9.590 2.100 11.340 2.260 ;
        RECT  12.060 1.340 12.300 1.620 ;
        RECT  12.100 1.340 12.300 2.000 ;
        RECT  11.180 1.840 12.300 2.000 ;
        RECT  2.760 0.440 3.950 0.600 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 0.900 1.020 1.100 ;
        RECT  0.100 2.100 1.020 2.300 ;
        RECT  0.100 0.900 0.300 2.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.280 1.460 8.700 1.680 ;
        RECT  8.280 1.520 10.000 1.680 ;
        RECT  9.840 1.680 11.000 1.840 ;
        RECT  8.500 1.140 8.700 1.680 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.960 1.200 11.340 1.360 ;
        RECT  11.180 1.200 11.340 1.560 ;
        RECT  11.180 1.400 11.640 1.560 ;
        RECT  9.700 0.790 9.900 1.360 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.580 0.400 ;
        RECT  4.210 -0.280 4.490 0.400 ;
        RECT  5.660 -0.280 5.940 0.400 ;
        RECT  8.520 -0.280 8.680 0.460 ;
        RECT  9.500 -0.280 9.780 0.400 ;
        RECT  10.620 -0.280 10.900 0.400 ;
        RECT  12.540 -0.280 12.820 0.400 ;
        RECT  13.620 -0.280 13.900 0.580 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 2.800 1.580 3.480 ;
        RECT  4.210 2.800 4.490 3.480 ;
        RECT  5.260 2.740 5.420 3.480 ;
        RECT  9.020 2.740 9.780 3.480 ;
        RECT  10.620 2.800 10.900 3.480 ;
        RECT  12.540 2.800 12.820 3.480 ;
        RECT  13.620 2.620 13.900 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  11.500 2.160 12.940 2.320 ;
        RECT  12.780 0.880 12.940 2.320 ;
        RECT  11.540 0.880 12.940 1.040 ;
        RECT  10.060 0.560 12.340 0.720 ;
        RECT  10.060 2.480 12.340 2.640 ;
        RECT  5.900 2.280 8.500 2.440 ;
        RECT  8.340 2.000 8.500 2.440 ;
        RECT  7.380 1.960 7.700 2.440 ;
        RECT  5.900 1.250 6.060 2.440 ;
        RECT  8.340 2.000 9.300 2.160 ;
        RECT  7.380 0.440 7.540 2.440 ;
        RECT  5.900 1.250 6.220 1.530 ;
        RECT  8.200 0.730 9.300 0.890 ;
        RECT  8.200 0.440 8.360 0.890 ;
        RECT  7.380 0.440 8.360 0.600 ;
        RECT  7.880 1.840 8.180 2.060 ;
        RECT  7.880 0.760 8.040 2.060 ;
        RECT  7.820 1.320 8.040 1.600 ;
        RECT  6.820 1.960 7.100 2.120 ;
        RECT  6.940 0.560 7.100 2.120 ;
        RECT  5.580 0.560 5.740 1.650 ;
        RECT  6.740 0.560 7.100 1.040 ;
        RECT  5.580 0.560 7.100 0.720 ;
        RECT  6.220 1.840 6.540 2.060 ;
        RECT  6.380 0.880 6.540 2.060 ;
        RECT  6.180 0.880 6.540 1.040 ;
        RECT  2.670 2.480 4.990 2.640 ;
        RECT  4.830 0.880 4.990 2.640 ;
        RECT  2.670 1.080 2.830 2.640 ;
        RECT  4.030 1.380 4.990 1.540 ;
        RECT  2.450 1.080 2.830 1.300 ;
        RECT  3.710 0.880 3.870 2.320 ;
        RECT  3.190 0.760 3.350 2.320 ;
        RECT  1.180 0.560 1.340 1.660 ;
        RECT  2.390 0.760 3.350 0.920 ;
        RECT  2.390 0.560 2.550 0.920 ;
        RECT  1.180 0.560 2.550 0.720 ;
        RECT  1.920 2.000 2.220 2.280 ;
        RECT  2.060 1.020 2.220 2.280 ;
        RECT  1.860 1.020 2.220 1.180 ;
    END
END FA1HHD

MACRO FA1KHD
    CLASS CORE ;
    FOREIGN FA1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  15.700 0.900 15.900 2.300 ;
        RECT  14.020 2.100 15.900 2.300 ;
        RECT  14.020 0.900 15.900 1.100 ;
        END
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.710 0.560 6.340 0.720 ;
        RECT  6.180 0.560 6.340 2.280 ;
        RECT  6.180 2.120 6.660 2.280 ;
        RECT  6.500 2.120 6.660 2.760 ;
        RECT  9.580 2.360 9.740 2.760 ;
        RECT  6.500 2.600 9.740 2.760 ;
        RECT  10.510 2.100 10.670 2.520 ;
        RECT  9.580 2.360 10.670 2.520 ;
        RECT  12.100 1.840 12.260 2.260 ;
        RECT  10.510 2.100 12.260 2.260 ;
        RECT  12.900 1.340 13.140 2.000 ;
        RECT  12.100 1.840 13.140 2.000 ;
        RECT  3.630 0.440 4.870 0.600 ;
        END
    END CI
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 0.900 1.940 1.100 ;
        RECT  0.100 2.100 1.940 2.300 ;
        RECT  0.100 0.900 0.300 2.300 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.200 1.460 9.500 1.680 ;
        RECT  9.200 1.520 11.920 1.680 ;
        RECT  9.300 1.140 9.500 1.680 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.880 1.200 12.260 1.360 ;
        RECT  12.100 1.200 12.260 1.560 ;
        RECT  12.100 1.400 12.560 1.560 ;
        RECT  10.500 0.790 10.700 1.360 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  2.220 -0.280 2.500 0.400 ;
        RECT  5.130 -0.280 5.410 0.400 ;
        RECT  6.580 -0.280 6.860 0.400 ;
        RECT  9.440 -0.280 9.600 0.460 ;
        RECT  10.420 -0.280 10.700 0.400 ;
        RECT  11.540 -0.280 11.820 0.400 ;
        RECT  13.460 -0.280 13.740 0.400 ;
        RECT  14.540 -0.280 14.820 0.580 ;
        RECT  15.580 -0.280 15.860 0.580 ;
        RECT  0.000 -0.280 16.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.620 1.420 3.480 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  5.130 2.800 5.410 3.480 ;
        RECT  6.180 2.740 6.340 3.480 ;
        RECT  9.940 2.800 10.220 3.480 ;
        RECT  10.420 2.800 10.700 3.480 ;
        RECT  9.940 2.880 10.700 3.480 ;
        RECT  11.540 2.800 11.820 3.480 ;
        RECT  13.460 2.800 13.740 3.480 ;
        RECT  14.540 2.620 14.820 3.480 ;
        RECT  15.580 2.620 15.860 3.480 ;
        RECT  0.000 2.920 16.000 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  12.420 2.160 13.860 2.320 ;
        RECT  13.700 0.880 13.860 2.320 ;
        RECT  12.460 0.880 13.860 1.040 ;
        RECT  10.980 0.560 13.260 0.720 ;
        RECT  10.980 2.480 13.260 2.640 ;
        RECT  6.820 2.280 9.420 2.440 ;
        RECT  9.260 2.000 9.420 2.440 ;
        RECT  8.300 1.960 8.620 2.440 ;
        RECT  6.820 1.400 6.980 2.440 ;
        RECT  9.260 2.000 10.220 2.160 ;
        RECT  8.300 0.440 8.460 2.440 ;
        RECT  6.820 1.400 7.140 1.680 ;
        RECT  9.120 0.730 10.220 0.890 ;
        RECT  9.120 0.440 9.280 0.890 ;
        RECT  8.300 0.440 9.280 0.600 ;
        RECT  8.800 1.840 9.100 2.060 ;
        RECT  8.800 0.760 8.960 2.060 ;
        RECT  8.740 1.320 8.960 1.600 ;
        RECT  7.740 1.960 8.020 2.120 ;
        RECT  7.860 0.560 8.020 2.120 ;
        RECT  6.500 0.560 6.660 1.650 ;
        RECT  7.660 0.560 8.020 1.040 ;
        RECT  6.500 0.560 8.020 0.720 ;
        RECT  7.140 1.840 7.460 2.060 ;
        RECT  7.300 0.880 7.460 2.060 ;
        RECT  7.100 0.880 7.460 1.040 ;
        RECT  3.590 2.480 5.910 2.640 ;
        RECT  5.750 0.880 5.910 2.640 ;
        RECT  3.590 1.080 3.750 2.640 ;
        RECT  4.970 1.430 5.250 1.650 ;
        RECT  4.970 1.430 5.910 1.590 ;
        RECT  3.370 1.080 3.750 1.300 ;
        RECT  4.630 0.880 4.790 2.320 ;
        RECT  4.110 0.760 4.270 2.320 ;
        RECT  2.100 0.560 2.260 1.670 ;
        RECT  3.310 0.760 4.270 0.920 ;
        RECT  3.310 0.560 3.470 0.920 ;
        RECT  2.100 0.560 3.470 0.720 ;
        RECT  2.840 2.040 3.140 2.320 ;
        RECT  2.980 1.020 3.140 2.320 ;
        RECT  2.780 1.020 3.140 1.180 ;
    END
END FA1KHD

MACRO FILLER16EHD
    CLASS CORE SPACER ;
    FOREIGN FILLER16EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  5.620 -0.280 6.280 0.400 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  6.020 2.800 6.300 3.480 ;
        RECT  0.120 2.800 0.780 3.480 ;
        END
    END VCC
END FILLER16EHD

MACRO FILLER1HD
    CLASS CORE SPACER ;
    FOREIGN FILLER1HD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 0.400 0.280 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 0.400 3.480 ;
        END
    END VCC
END FILLER1HD

MACRO FILLER2HD
    CLASS CORE SPACER ;
    FOREIGN FILLER2HD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 0.800 0.280 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 0.800 3.480 ;
        END
    END VCC
END FILLER2HD

MACRO FILLER32EHD
    CLASS CORE SPACER ;
    FOREIGN FILLER32EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        RECT  12.420 -0.280 12.700 0.400 ;
        RECT  5.880 -0.280 6.920 0.400 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 12.800 3.480 ;
        RECT  12.020 2.800 12.680 3.480 ;
        RECT  6.260 2.800 6.540 3.480 ;
        RECT  0.120 2.800 0.780 3.480 ;
        END
    END VCC
END FILLER32EHD

MACRO FILLER3HD
    CLASS CORE SPACER ;
    FOREIGN FILLER3HD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        END
    END VCC
END FILLER3HD

MACRO FILLER4EHD
    CLASS CORE SPACER ;
    FOREIGN FILLER4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 1.480 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.120 2.800 1.500 3.480 ;
        END
    END VCC
END FILLER4EHD

MACRO FILLER64EHD
    CLASS CORE SPACER ;
    FOREIGN FILLER64EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 25.600 0.280 ;
        RECT  25.220 -0.280 25.500 0.400 ;
        RECT  18.550 -0.280 19.590 0.400 ;
        RECT  12.660 -0.280 12.940 0.400 ;
        RECT  6.010 -0.280 7.050 0.400 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 25.600 3.480 ;
        RECT  24.820 2.800 25.480 3.480 ;
        RECT  18.930 2.800 19.210 3.480 ;
        RECT  12.280 2.800 13.320 3.480 ;
        RECT  6.390 2.800 6.670 3.480 ;
        RECT  0.120 2.800 0.780 3.480 ;
        END
    END VCC
END FILLER64EHD

MACRO FILLER8EHD
    CLASS CORE SPACER ;
    FOREIGN FILLER8EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  2.420 -0.280 3.080 0.400 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  2.820 2.800 3.100 3.480 ;
        RECT  0.120 2.800 0.780 3.480 ;
        END
    END VCC
END FILLER8EHD

MACRO GCBETCHD
    CLASS CORE ;
    FOREIGN GCBETCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.470 1.430 6.700 1.710 ;
        RECT  6.500 1.030 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.270 2.000 1.550 ;
        RECT  1.700 0.920 1.900 1.880 ;
        END
    END E
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.860 7.500 2.460 ;
        RECT  5.630 2.300 7.500 2.460 ;
        RECT  7.280 0.860 7.500 1.140 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.620 -0.280 1.900 0.400 ;
        RECT  3.820 -0.280 4.100 0.600 ;
        RECT  6.140 -0.280 6.420 0.480 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 2.730 4.540 3.480 ;
        RECT  6.550 2.620 6.830 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.620 2.620 1.750 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.420 1.980 7.110 2.140 ;
        RECT  6.950 1.430 7.110 2.140 ;
        RECT  5.420 1.340 5.580 2.140 ;
        RECT  5.570 0.640 6.980 0.800 ;
        RECT  5.100 0.440 5.260 2.530 ;
        RECT  5.900 0.960 6.060 1.620 ;
        RECT  5.100 0.960 6.060 1.120 ;
        RECT  3.640 0.820 4.420 0.980 ;
        RECT  4.260 0.440 4.420 0.980 ;
        RECT  4.260 0.440 5.260 0.600 ;
        RECT  1.910 2.600 4.160 2.760 ;
        RECT  4.000 2.410 4.160 2.760 ;
        RECT  1.910 2.300 2.070 2.760 ;
        RECT  4.000 2.410 4.940 2.570 ;
        RECT  4.780 1.340 4.940 2.570 ;
        RECT  0.100 2.300 2.070 2.460 ;
        RECT  0.820 0.920 0.980 2.460 ;
        RECT  3.440 1.340 4.940 1.500 ;
        RECT  0.160 0.920 0.980 1.080 ;
        RECT  0.160 0.540 0.320 1.080 ;
        RECT  2.800 2.280 3.840 2.440 ;
        RECT  3.680 1.890 3.840 2.440 ;
        RECT  2.800 0.760 2.960 2.440 ;
        RECT  3.680 1.890 4.620 2.050 ;
        RECT  2.760 0.760 2.960 1.040 ;
        RECT  3.120 1.840 3.520 2.120 ;
        RECT  3.120 0.440 3.280 2.120 ;
        RECT  3.120 0.440 3.620 0.600 ;
        RECT  1.200 1.840 1.400 2.120 ;
        RECT  1.200 0.560 1.360 2.120 ;
        RECT  1.200 0.560 2.600 0.720 ;
        RECT  2.440 0.440 2.840 0.600 ;
        RECT  2.240 0.880 2.400 2.260 ;
        RECT  2.180 0.880 2.460 1.040 ;
    END
END GCBETCHD

MACRO GCBETEHD
    CLASS CORE ;
    FOREIGN GCBETEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.470 1.430 6.700 1.710 ;
        RECT  6.500 1.030 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.270 2.000 1.550 ;
        RECT  1.700 0.920 1.900 1.880 ;
        END
    END E
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.880 9.100 2.340 ;
        RECT  8.880 2.060 9.100 2.340 ;
        RECT  8.860 0.880 9.100 1.160 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.620 -0.280 1.900 0.400 ;
        RECT  3.820 -0.280 4.100 0.600 ;
        RECT  6.140 -0.280 6.420 0.480 ;
        RECT  8.280 -0.280 8.560 1.060 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 2.730 4.540 3.480 ;
        RECT  6.550 2.620 6.830 3.480 ;
        RECT  8.300 2.620 8.580 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.620 2.620 1.750 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.770 1.860 7.960 2.140 ;
        RECT  7.800 0.880 7.960 2.140 ;
        RECT  8.460 1.420 8.740 1.640 ;
        RECT  7.800 1.420 8.740 1.580 ;
        RECT  5.630 2.300 7.500 2.460 ;
        RECT  7.300 0.860 7.500 2.460 ;
        RECT  7.300 1.430 7.590 1.710 ;
        RECT  7.280 0.860 7.500 1.140 ;
        RECT  5.420 1.980 7.110 2.140 ;
        RECT  6.950 1.430 7.110 2.140 ;
        RECT  5.420 1.340 5.580 2.140 ;
        RECT  5.570 0.640 6.980 0.800 ;
        RECT  5.100 0.440 5.260 2.530 ;
        RECT  5.900 0.960 6.060 1.620 ;
        RECT  5.100 0.960 6.060 1.120 ;
        RECT  3.640 0.820 4.420 0.980 ;
        RECT  4.260 0.440 4.420 0.980 ;
        RECT  4.260 0.440 5.260 0.600 ;
        RECT  1.910 2.600 4.160 2.760 ;
        RECT  4.000 2.410 4.160 2.760 ;
        RECT  1.910 2.300 2.070 2.760 ;
        RECT  4.000 2.410 4.940 2.570 ;
        RECT  4.780 1.340 4.940 2.570 ;
        RECT  0.100 2.300 2.070 2.460 ;
        RECT  0.820 0.920 0.980 2.460 ;
        RECT  3.440 1.340 4.940 1.500 ;
        RECT  0.160 0.920 0.980 1.080 ;
        RECT  0.160 0.540 0.320 1.080 ;
        RECT  2.800 2.280 3.840 2.440 ;
        RECT  3.680 1.890 3.840 2.440 ;
        RECT  2.800 0.760 2.960 2.440 ;
        RECT  3.680 1.890 4.620 2.050 ;
        RECT  2.760 0.760 2.960 1.040 ;
        RECT  3.120 1.840 3.520 2.120 ;
        RECT  3.120 0.440 3.280 2.120 ;
        RECT  3.120 0.440 3.620 0.600 ;
        RECT  1.200 1.840 1.400 2.120 ;
        RECT  1.200 0.560 1.360 2.120 ;
        RECT  1.200 0.560 2.600 0.720 ;
        RECT  2.440 0.440 2.840 0.600 ;
        RECT  2.240 0.880 2.400 2.260 ;
        RECT  2.180 0.880 2.460 1.040 ;
    END
END GCBETEHD

MACRO GCBETHHD
    CLASS CORE ;
    FOREIGN GCBETHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.410 1.430 6.700 1.710 ;
        RECT  6.500 1.030 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.270 2.000 1.550 ;
        RECT  1.700 0.920 1.900 1.880 ;
        END
    END E
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.880 9.100 2.340 ;
        RECT  8.760 2.060 9.100 2.340 ;
        RECT  8.760 0.880 9.100 1.160 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.620 -0.280 1.900 0.400 ;
        RECT  3.820 -0.280 4.100 0.600 ;
        RECT  6.080 -0.280 6.360 0.480 ;
        RECT  8.180 -0.280 8.460 1.060 ;
        RECT  9.280 -0.280 9.440 1.040 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 2.730 4.540 3.480 ;
        RECT  6.490 2.620 6.770 3.480 ;
        RECT  8.180 2.620 8.460 3.480 ;
        RECT  9.220 2.620 9.500 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.620 2.620 1.750 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.670 2.050 7.860 2.330 ;
        RECT  7.700 0.880 7.860 2.330 ;
        RECT  7.700 1.420 8.640 1.580 ;
        RECT  5.570 2.300 7.510 2.460 ;
        RECT  7.350 0.860 7.510 2.460 ;
        RECT  7.310 1.430 7.530 1.710 ;
        RECT  7.220 0.860 7.510 1.140 ;
        RECT  5.360 1.980 7.050 2.140 ;
        RECT  6.890 1.430 7.050 2.140 ;
        RECT  5.360 1.310 5.520 2.140 ;
        RECT  5.510 0.640 6.920 0.800 ;
        RECT  5.040 0.440 5.200 2.530 ;
        RECT  5.840 0.960 6.000 1.620 ;
        RECT  5.040 0.960 6.000 1.120 ;
        RECT  3.640 0.820 4.420 0.980 ;
        RECT  4.260 0.440 4.420 0.980 ;
        RECT  4.260 0.440 5.200 0.600 ;
        RECT  1.910 2.600 4.160 2.760 ;
        RECT  4.000 2.410 4.160 2.760 ;
        RECT  1.910 2.300 2.070 2.760 ;
        RECT  4.000 2.410 4.880 2.570 ;
        RECT  4.720 1.250 4.880 2.570 ;
        RECT  0.100 2.300 2.070 2.460 ;
        RECT  0.820 0.920 0.980 2.460 ;
        RECT  3.440 1.300 4.880 1.460 ;
        RECT  4.600 1.250 4.880 1.460 ;
        RECT  0.160 0.920 0.980 1.080 ;
        RECT  0.160 0.540 0.320 1.080 ;
        RECT  2.800 2.280 3.840 2.440 ;
        RECT  3.680 1.850 3.840 2.440 ;
        RECT  2.800 0.760 2.960 2.440 ;
        RECT  3.680 1.850 4.560 2.010 ;
        RECT  4.340 1.680 4.560 2.010 ;
        RECT  2.760 0.760 2.960 1.040 ;
        RECT  3.120 1.840 3.520 2.120 ;
        RECT  3.120 0.440 3.280 2.120 ;
        RECT  3.120 0.440 3.620 0.600 ;
        RECT  1.200 1.840 1.400 2.120 ;
        RECT  1.200 0.560 1.360 2.120 ;
        RECT  1.200 0.560 2.600 0.720 ;
        RECT  2.440 0.440 2.840 0.600 ;
        RECT  2.240 0.880 2.400 2.260 ;
        RECT  2.180 0.880 2.460 1.040 ;
    END
END GCBETHHD

MACRO GCBETKHD
    CLASS CORE ;
    FOREIGN GCBETKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.410 1.430 6.700 1.710 ;
        RECT  6.500 1.030 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.270 2.000 1.550 ;
        RECT  1.700 0.920 1.900 1.880 ;
        END
    END E
    PIN CKB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END CKB
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.800 0.880 8.960 2.280 ;
        RECT  9.700 0.880 9.900 2.280 ;
        RECT  9.700 0.880 9.960 1.160 ;
        RECT  8.700 2.120 10.060 2.280 ;
        RECT  8.760 0.880 8.960 1.160 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.620 -0.280 1.900 0.400 ;
        RECT  3.820 -0.280 4.100 0.600 ;
        RECT  6.080 -0.280 6.360 0.480 ;
        RECT  8.180 -0.280 8.460 1.060 ;
        RECT  9.280 -0.280 9.440 1.000 ;
        RECT  10.320 -0.280 10.480 1.000 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.320 2.730 4.540 3.480 ;
        RECT  6.490 2.620 6.770 3.480 ;
        RECT  8.180 2.620 8.460 3.480 ;
        RECT  9.220 2.620 9.500 3.480 ;
        RECT  10.260 2.620 10.540 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.620 2.620 1.750 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.670 2.050 7.860 2.330 ;
        RECT  7.700 0.880 7.860 2.330 ;
        RECT  7.700 1.420 8.640 1.580 ;
        RECT  5.570 2.300 7.510 2.460 ;
        RECT  7.350 0.860 7.510 2.460 ;
        RECT  7.310 1.430 7.530 1.710 ;
        RECT  7.220 0.860 7.510 1.140 ;
        RECT  5.360 1.980 7.050 2.140 ;
        RECT  6.890 1.430 7.050 2.140 ;
        RECT  5.360 1.310 5.520 2.140 ;
        RECT  5.510 0.640 6.920 0.800 ;
        RECT  5.040 0.440 5.200 2.530 ;
        RECT  5.840 0.960 6.000 1.620 ;
        RECT  5.040 0.960 6.000 1.120 ;
        RECT  3.640 0.820 4.420 0.980 ;
        RECT  4.260 0.440 4.420 0.980 ;
        RECT  4.260 0.440 5.200 0.600 ;
        RECT  1.910 2.600 4.160 2.760 ;
        RECT  4.000 2.410 4.160 2.760 ;
        RECT  1.910 2.300 2.070 2.760 ;
        RECT  4.000 2.410 4.880 2.570 ;
        RECT  4.720 1.250 4.880 2.570 ;
        RECT  0.100 2.300 2.070 2.460 ;
        RECT  0.820 0.920 0.980 2.460 ;
        RECT  3.440 1.300 4.880 1.460 ;
        RECT  4.600 1.250 4.880 1.460 ;
        RECT  0.160 0.920 0.980 1.080 ;
        RECT  0.160 0.540 0.320 1.080 ;
        RECT  2.800 2.280 3.840 2.440 ;
        RECT  3.680 1.850 3.840 2.440 ;
        RECT  2.800 0.760 2.960 2.440 ;
        RECT  3.680 1.850 4.560 2.010 ;
        RECT  4.340 1.680 4.560 2.010 ;
        RECT  2.760 0.760 2.960 1.040 ;
        RECT  3.120 1.840 3.520 2.120 ;
        RECT  3.120 0.440 3.280 2.120 ;
        RECT  3.120 0.440 3.630 0.600 ;
        RECT  1.200 1.840 1.400 2.120 ;
        RECT  1.200 0.560 1.360 2.120 ;
        RECT  1.200 0.560 2.600 0.720 ;
        RECT  2.440 0.440 2.840 0.600 ;
        RECT  2.240 0.880 2.400 2.260 ;
        RECT  2.180 0.880 2.460 1.040 ;
    END
END GCBETKHD

MACRO GCKETCHD
    CLASS CORE ;
    FOREIGN GCKETCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.880 1.340 5.100 1.620 ;
        RECT  4.900 0.960 7.060 1.120 ;
        RECT  6.900 0.960 7.060 1.750 ;
        RECT  4.900 0.960 5.100 1.620 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.430 6.700 1.960 ;
        RECT  6.420 1.430 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.270 0.440 1.550 ;
        RECT  0.100 0.920 0.300 1.880 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.640 2.060 7.900 2.340 ;
        RECT  7.700 0.860 7.930 1.140 ;
        RECT  7.700 0.860 7.900 2.340 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 -0.280 2.660 0.400 ;
        RECT  4.490 -0.280 4.770 0.400 ;
        RECT  6.100 -0.280 6.380 0.480 ;
        RECT  8.230 -0.280 8.510 1.020 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.800 2.730 3.020 3.480 ;
        RECT  4.000 2.800 4.800 3.480 ;
        RECT  6.560 2.620 6.840 3.480 ;
        RECT  8.100 2.220 8.380 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.740 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.640 2.600 6.400 2.760 ;
        RECT  6.240 2.300 6.400 2.760 ;
        RECT  6.240 2.300 7.440 2.460 ;
        RECT  7.280 0.860 7.440 2.460 ;
        RECT  7.280 1.340 7.540 1.620 ;
        RECT  7.280 0.860 7.450 1.140 ;
        RECT  5.530 0.640 6.940 0.800 ;
        RECT  3.580 0.920 3.740 2.490 ;
        RECT  3.580 2.280 5.720 2.440 ;
        RECT  5.560 1.460 5.720 2.440 ;
        RECT  5.560 1.460 6.070 1.620 ;
        RECT  5.910 1.340 6.070 1.620 ;
        RECT  3.000 0.920 3.280 1.120 ;
        RECT  2.220 0.920 3.740 1.080 ;
        RECT  4.480 1.900 5.400 2.060 ;
        RECT  4.480 0.560 4.640 2.060 ;
        RECT  4.400 1.440 4.640 1.720 ;
        RECT  5.050 0.560 5.330 0.760 ;
        RECT  1.650 0.560 5.330 0.720 ;
        RECT  1.000 0.440 1.810 0.600 ;
        RECT  3.950 1.840 4.220 2.120 ;
        RECT  3.950 0.940 4.110 2.120 ;
        RECT  3.900 1.380 4.110 1.660 ;
        RECT  1.000 2.600 2.640 2.760 ;
        RECT  2.480 2.410 2.640 2.760 ;
        RECT  2.480 2.410 3.420 2.570 ;
        RECT  3.260 1.340 3.420 2.570 ;
        RECT  1.920 1.460 3.420 1.620 ;
        RECT  3.140 1.340 3.420 1.620 ;
        RECT  1.280 2.280 2.320 2.440 ;
        RECT  2.160 1.890 2.320 2.440 ;
        RECT  1.280 0.820 1.440 2.440 ;
        RECT  2.160 1.890 3.100 2.050 ;
        RECT  1.600 1.840 2.000 2.120 ;
        RECT  1.600 0.880 1.760 2.120 ;
        RECT  1.600 0.880 2.060 1.040 ;
        RECT  0.720 0.880 0.880 2.260 ;
        RECT  0.660 0.880 0.940 1.040 ;
    END
END GCKETCHD

MACRO GCKETEHD
    CLASS CORE ;
    FOREIGN GCKETEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.880 1.340 5.100 1.620 ;
        RECT  4.900 0.960 7.060 1.120 ;
        RECT  6.900 0.960 7.060 1.750 ;
        RECT  4.900 0.960 5.100 1.620 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.430 6.700 1.960 ;
        RECT  6.420 1.430 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.270 0.440 1.550 ;
        RECT  0.100 0.920 0.300 1.880 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.640 2.060 7.900 2.340 ;
        RECT  7.700 0.860 7.930 1.140 ;
        RECT  7.700 0.860 7.900 2.340 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 -0.280 2.660 0.400 ;
        RECT  4.490 -0.280 4.770 0.400 ;
        RECT  6.100 -0.280 6.380 0.480 ;
        RECT  8.230 -0.280 8.510 1.020 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.800 2.730 3.020 3.480 ;
        RECT  4.000 2.800 4.800 3.480 ;
        RECT  6.560 2.620 6.840 3.480 ;
        RECT  8.100 2.620 8.380 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.740 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.640 2.600 6.400 2.760 ;
        RECT  6.240 2.300 6.400 2.760 ;
        RECT  6.240 2.300 7.440 2.460 ;
        RECT  7.280 0.860 7.440 2.460 ;
        RECT  7.280 1.340 7.540 1.620 ;
        RECT  7.280 0.860 7.450 1.140 ;
        RECT  5.530 0.640 6.940 0.800 ;
        RECT  3.580 0.920 3.740 2.490 ;
        RECT  3.580 2.280 5.720 2.440 ;
        RECT  5.560 1.460 5.720 2.440 ;
        RECT  5.560 1.460 6.070 1.620 ;
        RECT  5.910 1.340 6.070 1.620 ;
        RECT  3.000 0.920 3.280 1.120 ;
        RECT  2.220 0.920 3.740 1.080 ;
        RECT  4.480 1.900 5.400 2.060 ;
        RECT  4.480 0.560 4.640 2.060 ;
        RECT  4.400 1.440 4.640 1.720 ;
        RECT  5.050 0.560 5.330 0.760 ;
        RECT  1.650 0.560 5.330 0.720 ;
        RECT  1.000 0.440 1.810 0.600 ;
        RECT  3.950 1.840 4.220 2.120 ;
        RECT  3.950 0.940 4.110 2.120 ;
        RECT  3.900 1.380 4.110 1.660 ;
        RECT  1.000 2.600 2.640 2.760 ;
        RECT  2.480 2.410 2.640 2.760 ;
        RECT  2.480 2.410 3.420 2.570 ;
        RECT  3.260 1.340 3.420 2.570 ;
        RECT  1.920 1.460 3.420 1.620 ;
        RECT  3.140 1.340 3.420 1.620 ;
        RECT  1.280 2.280 2.320 2.440 ;
        RECT  2.160 1.890 2.320 2.440 ;
        RECT  1.280 0.820 1.440 2.440 ;
        RECT  2.160 1.890 3.100 2.050 ;
        RECT  1.600 1.840 2.000 2.120 ;
        RECT  1.600 0.880 1.760 2.120 ;
        RECT  1.600 0.880 2.060 1.040 ;
        RECT  0.720 0.880 0.880 2.260 ;
        RECT  0.660 0.880 0.940 1.040 ;
    END
END GCKETEHD

MACRO GCKETHHD
    CLASS CORE ;
    FOREIGN GCKETHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.880 1.340 5.100 1.620 ;
        RECT  4.900 0.960 7.060 1.120 ;
        RECT  6.900 0.960 7.060 1.750 ;
        RECT  4.900 0.960 5.100 1.620 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.430 6.700 1.960 ;
        RECT  6.420 1.430 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.270 0.440 1.550 ;
        RECT  0.100 0.920 0.300 1.880 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.640 2.060 7.880 2.340 ;
        RECT  7.720 0.860 7.930 1.140 ;
        RECT  8.810 0.860 9.100 1.140 ;
        RECT  8.900 0.860 9.100 2.280 ;
        RECT  7.640 2.120 9.100 2.280 ;
        RECT  7.720 0.860 7.880 2.340 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 -0.280 2.660 0.400 ;
        RECT  4.490 -0.280 4.770 0.400 ;
        RECT  6.100 -0.280 6.380 0.480 ;
        RECT  8.230 -0.280 8.510 1.020 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.800 2.730 3.020 3.480 ;
        RECT  4.000 2.800 4.800 3.480 ;
        RECT  6.560 2.620 6.840 3.480 ;
        RECT  8.100 2.620 8.380 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  0.100 2.740 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.640 2.600 6.400 2.760 ;
        RECT  6.240 2.300 6.400 2.760 ;
        RECT  6.240 2.300 7.440 2.460 ;
        RECT  7.280 0.860 7.440 2.460 ;
        RECT  7.280 1.340 7.540 1.620 ;
        RECT  7.280 0.860 7.450 1.140 ;
        RECT  5.530 0.640 6.940 0.800 ;
        RECT  3.580 0.920 3.740 2.490 ;
        RECT  3.580 2.280 5.720 2.440 ;
        RECT  5.560 1.460 5.720 2.440 ;
        RECT  5.560 1.460 6.070 1.620 ;
        RECT  5.910 1.340 6.070 1.620 ;
        RECT  3.000 0.920 3.280 1.120 ;
        RECT  2.220 0.920 3.740 1.080 ;
        RECT  4.480 1.900 5.400 2.060 ;
        RECT  4.480 0.560 4.640 2.060 ;
        RECT  4.400 1.440 4.640 1.720 ;
        RECT  5.050 0.560 5.330 0.760 ;
        RECT  1.650 0.560 5.330 0.720 ;
        RECT  1.000 0.440 1.810 0.600 ;
        RECT  3.950 1.840 4.220 2.120 ;
        RECT  3.950 0.940 4.110 2.120 ;
        RECT  3.900 1.380 4.110 1.660 ;
        RECT  1.000 2.600 2.640 2.760 ;
        RECT  2.480 2.410 2.640 2.760 ;
        RECT  2.480 2.410 3.420 2.570 ;
        RECT  3.260 1.340 3.420 2.570 ;
        RECT  1.920 1.460 3.420 1.620 ;
        RECT  3.140 1.340 3.420 1.620 ;
        RECT  1.280 2.280 2.320 2.440 ;
        RECT  2.160 1.890 2.320 2.440 ;
        RECT  1.280 0.820 1.440 2.440 ;
        RECT  2.160 1.890 3.100 2.050 ;
        RECT  1.600 1.840 2.000 2.120 ;
        RECT  1.600 0.880 1.760 2.120 ;
        RECT  1.600 0.880 2.060 1.040 ;
        RECT  0.720 0.880 0.880 2.260 ;
        RECT  0.660 0.880 0.940 1.040 ;
    END
END GCKETHHD

MACRO GCKETKHD
    CLASS CORE ;
    FOREIGN GCKETKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.880 1.340 5.100 1.620 ;
        RECT  4.900 0.960 7.060 1.120 ;
        RECT  6.900 0.960 7.060 1.750 ;
        RECT  4.900 0.960 5.100 1.620 ;
        END
    END CK
    PIN TE
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.430 6.700 1.960 ;
        RECT  6.420 1.430 6.700 1.710 ;
        END
    END TE
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.270 0.440 1.550 ;
        RECT  0.100 0.920 0.300 1.880 ;
        END
    END E
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.580 2.060 7.880 2.280 ;
        RECT  7.720 0.860 7.930 1.140 ;
        RECT  8.810 0.860 9.100 1.140 ;
        RECT  8.900 0.860 9.100 2.280 ;
        RECT  9.720 0.860 9.880 2.280 ;
        RECT  7.580 2.120 9.980 2.280 ;
        RECT  9.720 0.860 10.010 1.140 ;
        RECT  7.720 0.860 7.880 2.280 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.380 -0.280 2.660 0.400 ;
        RECT  4.490 -0.280 4.770 0.400 ;
        RECT  6.100 -0.280 6.380 0.480 ;
        RECT  8.230 -0.280 8.510 1.020 ;
        RECT  9.270 -0.280 9.550 1.020 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.800 2.730 3.020 3.480 ;
        RECT  4.000 2.800 4.800 3.480 ;
        RECT  6.560 2.620 6.840 3.480 ;
        RECT  8.100 2.620 8.380 3.480 ;
        RECT  9.140 2.620 9.420 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.100 2.740 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.640 2.600 6.400 2.760 ;
        RECT  6.240 2.300 6.400 2.760 ;
        RECT  6.240 2.300 7.420 2.460 ;
        RECT  7.260 0.860 7.420 2.460 ;
        RECT  7.260 1.340 7.540 1.620 ;
        RECT  7.240 0.860 7.420 1.140 ;
        RECT  5.530 0.640 6.940 0.800 ;
        RECT  3.580 0.920 3.740 2.490 ;
        RECT  3.580 2.280 5.720 2.440 ;
        RECT  5.560 1.460 5.720 2.440 ;
        RECT  5.560 1.460 6.070 1.620 ;
        RECT  5.910 1.340 6.070 1.620 ;
        RECT  3.000 0.920 3.280 1.120 ;
        RECT  2.220 0.920 3.740 1.080 ;
        RECT  4.480 1.900 5.400 2.060 ;
        RECT  4.480 0.560 4.640 2.060 ;
        RECT  4.400 1.440 4.640 1.720 ;
        RECT  5.050 0.560 5.330 0.760 ;
        RECT  1.650 0.560 5.330 0.720 ;
        RECT  1.000 0.440 1.810 0.600 ;
        RECT  3.950 1.840 4.220 2.120 ;
        RECT  3.950 0.940 4.110 2.120 ;
        RECT  3.900 1.380 4.110 1.660 ;
        RECT  1.000 2.600 2.640 2.760 ;
        RECT  2.480 2.410 2.640 2.760 ;
        RECT  2.480 2.410 3.420 2.570 ;
        RECT  3.260 1.340 3.420 2.570 ;
        RECT  1.920 1.460 3.420 1.620 ;
        RECT  3.140 1.340 3.420 1.620 ;
        RECT  1.280 2.280 2.320 2.440 ;
        RECT  2.160 1.890 2.320 2.440 ;
        RECT  1.280 0.820 1.440 2.440 ;
        RECT  2.160 1.890 3.100 2.050 ;
        RECT  1.600 1.840 2.000 2.120 ;
        RECT  1.600 0.880 1.760 2.120 ;
        RECT  1.600 0.880 2.060 1.040 ;
        RECT  0.720 0.880 0.880 2.260 ;
        RECT  0.660 0.880 0.940 1.040 ;
    END
END GCKETKHD

MACRO HA1CHD
    CLASS CORE ;
    FOREIGN HA1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.780 0.620 5.500 0.820 ;
        RECT  5.300 0.620 5.500 2.040 ;
        RECT  4.960 1.840 5.500 2.040 ;
        RECT  4.960 1.840 5.180 2.120 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.650 6.300 2.440 ;
        RECT  6.080 2.160 6.300 2.440 ;
        RECT  6.080 0.650 6.300 0.930 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.220 0.700 1.840 ;
        RECT  0.520 1.060 1.260 1.220 ;
        RECT  1.100 0.440 1.260 1.220 ;
        RECT  1.100 0.440 2.740 0.600 ;
        RECT  2.580 0.570 3.330 0.730 ;
        RECT  3.170 0.570 3.330 1.680 ;
        RECT  3.170 1.520 4.310 1.680 ;
        RECT  0.480 1.410 0.700 1.690 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.410 1.500 1.960 ;
        RECT  1.280 1.410 1.500 1.690 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.510 -0.280 3.670 1.000 ;
        RECT  5.400 -0.280 5.680 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.340 2.800 3.620 3.480 ;
        RECT  4.340 2.620 4.620 3.480 ;
        RECT  5.460 2.740 5.740 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.860 1.900 1.140 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.300 2.280 5.890 2.440 ;
        RECT  5.730 1.370 5.890 2.440 ;
        RECT  2.300 0.970 2.460 2.440 ;
        RECT  2.240 0.970 2.520 1.130 ;
        RECT  3.740 1.900 4.730 2.060 ;
        RECT  4.570 1.020 4.730 2.060 ;
        RECT  4.360 1.020 4.730 1.180 ;
        RECT  4.360 0.680 4.520 1.180 ;
        RECT  1.660 2.600 3.180 2.760 ;
        RECT  1.660 0.960 1.820 2.760 ;
        RECT  2.820 0.910 2.980 2.120 ;
        RECT  0.100 2.540 0.380 2.760 ;
        RECT  0.160 0.600 0.320 2.760 ;
    END
END HA1CHD

MACRO HA1EHD
    CLASS CORE ;
    FOREIGN HA1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.040 1.840 5.260 2.120 ;
        RECT  5.040 0.940 5.500 1.140 ;
        RECT  5.300 0.940 5.500 2.040 ;
        RECT  5.040 1.840 5.500 2.040 ;
        RECT  5.040 0.860 5.200 1.140 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.650 6.300 2.450 ;
        RECT  6.080 2.170 6.300 2.450 ;
        RECT  6.080 0.650 6.300 0.930 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.220 0.700 1.840 ;
        RECT  0.520 1.060 1.260 1.220 ;
        RECT  1.100 0.440 1.260 1.220 ;
        RECT  1.100 0.440 2.740 0.600 ;
        RECT  2.580 0.570 3.330 0.730 ;
        RECT  3.170 0.570 3.330 1.680 ;
        RECT  3.170 1.520 4.400 1.680 ;
        RECT  0.480 1.410 0.700 1.690 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.410 1.500 1.960 ;
        RECT  1.280 1.410 1.500 1.690 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.510 -0.280 3.670 0.970 ;
        RECT  5.500 -0.280 5.780 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.340 2.800 3.620 3.480 ;
        RECT  4.340 2.620 4.620 3.480 ;
        RECT  5.500 2.620 5.780 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.860 1.940 1.140 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.300 2.280 5.890 2.440 ;
        RECT  5.730 1.370 5.890 2.440 ;
        RECT  2.300 0.970 2.460 2.440 ;
        RECT  5.680 1.370 5.900 1.690 ;
        RECT  2.240 0.970 2.520 1.130 ;
        RECT  3.740 1.900 4.880 2.060 ;
        RECT  4.720 1.020 4.880 2.060 ;
        RECT  4.460 1.020 4.880 1.180 ;
        RECT  1.660 2.600 3.180 2.760 ;
        RECT  1.660 0.960 1.820 2.760 ;
        RECT  2.820 0.910 2.980 2.120 ;
        RECT  0.100 2.540 0.380 2.760 ;
        RECT  0.160 0.600 0.320 2.760 ;
    END
END HA1EHD

MACRO HA1HHD
    CLASS CORE ;
    FOREIGN HA1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.860 6.300 2.120 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.900 7.500 2.300 ;
        RECT  7.100 2.100 7.500 2.300 ;
        RECT  7.100 0.900 7.500 1.100 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.140 0.700 1.840 ;
        RECT  1.570 1.140 1.850 1.560 ;
        RECT  1.860 0.520 2.020 1.300 ;
        RECT  0.500 1.140 2.020 1.300 ;
        RECT  1.860 0.520 3.730 0.680 ;
        RECT  3.570 0.520 3.730 1.680 ;
        RECT  3.570 1.520 5.440 1.680 ;
        RECT  0.480 1.410 0.700 1.690 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.170 1.740 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.910 -0.280 4.070 0.970 ;
        RECT  5.540 -0.280 5.820 0.580 ;
        RECT  6.580 -0.280 6.860 0.580 ;
        RECT  7.620 -0.280 7.900 0.580 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.080 2.600 4.240 3.480 ;
        RECT  5.540 2.620 5.820 3.480 ;
        RECT  6.580 2.620 6.860 3.480 ;
        RECT  7.620 2.620 7.900 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.670 2.420 0.950 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.720 2.280 6.840 2.440 ;
        RECT  6.680 1.470 6.840 2.440 ;
        RECT  1.710 2.280 3.600 2.440 ;
        RECT  3.440 1.840 3.600 2.440 ;
        RECT  4.720 1.840 4.880 2.440 ;
        RECT  2.750 0.960 2.910 2.440 ;
        RECT  1.710 2.220 1.990 2.440 ;
        RECT  3.440 1.840 4.880 2.000 ;
        RECT  6.680 1.470 7.090 1.630 ;
        RECT  2.700 0.960 2.910 1.240 ;
        RECT  5.040 1.840 5.260 2.120 ;
        RECT  5.040 1.900 5.940 2.060 ;
        RECT  5.780 1.020 5.940 2.060 ;
        RECT  4.900 1.020 5.940 1.180 ;
        RECT  4.400 2.600 4.840 2.760 ;
        RECT  2.500 2.600 3.920 2.760 ;
        RECT  3.760 2.160 3.920 2.760 ;
        RECT  4.400 2.160 4.560 2.760 ;
        RECT  3.760 2.160 4.560 2.320 ;
        RECT  3.070 1.840 3.280 2.120 ;
        RECT  3.070 0.960 3.230 2.120 ;
        RECT  3.070 0.960 3.400 1.240 ;
        RECT  1.250 2.130 1.490 2.410 ;
        RECT  1.330 1.780 1.490 2.410 ;
        RECT  1.330 1.780 2.590 1.940 ;
        RECT  2.180 1.660 2.590 1.940 ;
        RECT  2.180 0.960 2.340 1.940 ;
        RECT  0.160 0.540 0.320 2.160 ;
        RECT  1.480 0.500 1.700 0.780 ;
        RECT  0.160 0.580 1.700 0.740 ;
    END
END HA1HHD

MACRO HA1KHD
    CLASS CORE ;
    FOREIGN HA1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.520 1.840 6.920 2.120 ;
        RECT  6.920 1.020 7.080 2.060 ;
        RECT  6.520 1.020 7.820 1.180 ;
        RECT  6.520 1.900 7.820 2.060 ;
        RECT  6.520 0.860 6.740 1.180 ;
        END
    END C
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.900 9.500 2.300 ;
        RECT  8.860 0.900 10.180 1.100 ;
        RECT  8.900 2.100 10.180 2.300 ;
        RECT  8.920 2.080 9.080 2.360 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.140 0.700 1.840 ;
        RECT  0.500 1.140 2.020 1.300 ;
        RECT  1.860 0.520 2.020 1.560 ;
        RECT  1.740 1.140 2.020 1.560 ;
        RECT  1.860 0.520 4.130 0.680 ;
        RECT  3.970 0.520 4.130 1.680 ;
        RECT  3.970 1.520 5.840 1.680 ;
        RECT  0.480 1.410 0.700 1.690 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.170 1.740 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.310 -0.280 4.470 0.970 ;
        RECT  5.940 -0.280 6.220 0.580 ;
        RECT  6.980 -0.280 7.260 0.580 ;
        RECT  8.020 -0.280 8.300 0.580 ;
        RECT  9.380 -0.280 9.660 0.580 ;
        RECT  10.420 -0.280 10.700 0.580 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.480 2.600 4.640 3.480 ;
        RECT  5.940 2.620 6.220 3.480 ;
        RECT  6.980 2.620 7.260 3.480 ;
        RECT  8.020 2.620 8.300 3.480 ;
        RECT  9.380 2.620 9.660 3.480 ;
        RECT  10.420 2.620 10.700 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.840 2.580 1.120 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.120 2.280 8.680 2.440 ;
        RECT  8.520 1.370 8.680 2.440 ;
        RECT  1.880 2.280 4.000 2.440 ;
        RECT  3.840 1.840 4.000 2.440 ;
        RECT  5.120 1.840 5.280 2.440 ;
        RECT  3.150 0.960 3.310 2.440 ;
        RECT  1.880 2.220 2.160 2.440 ;
        RECT  3.840 1.840 5.280 2.000 ;
        RECT  3.100 0.960 3.310 1.240 ;
        RECT  5.440 1.840 5.660 2.120 ;
        RECT  5.440 1.900 6.340 2.060 ;
        RECT  6.180 1.020 6.340 2.060 ;
        RECT  5.300 1.020 6.340 1.180 ;
        RECT  4.800 2.600 5.320 2.760 ;
        RECT  2.500 2.600 4.320 2.760 ;
        RECT  4.160 2.160 4.320 2.760 ;
        RECT  4.800 2.160 4.960 2.760 ;
        RECT  4.160 2.160 4.960 2.320 ;
        RECT  3.470 1.840 3.680 2.120 ;
        RECT  3.470 0.960 3.630 2.120 ;
        RECT  3.470 0.960 3.800 1.240 ;
        RECT  1.420 2.130 1.660 2.410 ;
        RECT  1.500 1.780 1.660 2.410 ;
        RECT  1.500 1.780 2.990 1.940 ;
        RECT  2.180 1.660 2.990 1.940 ;
        RECT  2.180 0.960 2.340 1.940 ;
        RECT  0.160 0.540 0.320 2.160 ;
        RECT  1.480 0.500 1.700 0.780 ;
        RECT  0.160 0.580 1.700 0.740 ;
    END
END HA1KHD

MACRO INVCHD
    CLASS CORE ;
    FOREIGN INVCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 0.660 0.320 0.940 ;
        RECT  0.100 2.080 0.320 2.360 ;
        RECT  0.100 0.660 0.300 2.360 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.880 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        RECT  0.620 2.140 0.900 3.480 ;
        END
    END VCC
END INVCHD

MACRO INVCKDHD
    CLASS CORE ;
    FOREIGN INVCKDHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 0.540 1.100 2.280 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.460 1.600 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
END INVCKDHD

MACRO INVCKGHD
    CLASS CORE ;
    FOREIGN INVCKGHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.900 1.500 2.160 ;
        RECT  0.700 1.960 1.500 2.160 ;
        RECT  0.660 0.900 1.500 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.420 1.600 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  1.220 -0.280 1.500 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 2.320 1.500 3.480 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
END INVCKGHD

MACRO INVCKHHD
    CLASS CORE ;
    FOREIGN INVCKHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.900 1.900 2.280 ;
        RECT  0.660 2.080 1.900 2.280 ;
        RECT  0.860 0.900 1.900 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.420 1.600 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.620 -0.280 1.900 0.400 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.260 2.440 1.900 3.480 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
END INVCKHHD

MACRO INVCKIHD
    CLASS CORE ;
    FOREIGN INVCKIHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.760 1.550 2.280 1.800 ;
        RECT  2.080 0.880 2.280 1.160 ;
        RECT  2.120 0.880 2.280 2.340 ;
        RECT  2.080 1.550 2.280 2.340 ;
        RECT  0.760 0.840 0.920 2.700 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.420 1.600 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.580 0.400 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 2.800 1.580 3.480 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
END INVCKIHD

MACRO INVCKJHD
    CLASS CORE ;
    FOREIGN INVCKJHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.760 1.500 2.680 1.800 ;
        RECT  2.480 0.880 2.680 2.320 ;
        RECT  0.760 0.800 0.920 2.480 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.380 0.460 1.540 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.270 -0.280 1.970 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.390 2.580 2.030 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
END INVCKJHD

MACRO INVCKKHD
    CLASS CORE ;
    FOREIGN INVCKKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.680 2.080 0.920 2.360 ;
        RECT  2.320 0.920 2.680 1.870 ;
        RECT  0.760 1.470 2.680 1.870 ;
        RECT  2.360 0.920 2.680 2.360 ;
        RECT  0.760 0.890 0.920 2.360 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.400 0.480 1.560 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.940 0.680 ;
        RECT  2.820 -0.280 3.100 0.690 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.280 2.580 1.920 3.480 ;
        RECT  2.820 2.620 3.100 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVCKKHD

MACRO INVCKLHD
    CLASS CORE ;
    FOREIGN INVCKLHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.880 0.830 1.040 2.360 ;
        RECT  0.680 2.080 1.040 2.360 ;
        RECT  2.260 0.790 2.420 2.360 ;
        RECT  2.240 1.290 2.420 2.360 ;
        RECT  0.880 1.290 3.480 1.890 ;
        RECT  3.280 0.790 3.480 2.360 ;
        RECT  0.720 0.830 1.040 1.110 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.680 1.620 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.900 0.680 ;
        RECT  2.760 -0.280 3.400 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.580 1.860 3.480 ;
        RECT  2.700 2.620 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVCKLHD

MACRO INVCKMHD
    CLASS CORE ;
    FOREIGN INVCKMHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.000 0.880 1.160 2.360 ;
        RECT  0.680 2.080 1.160 2.360 ;
        RECT  2.480 0.790 2.640 2.360 ;
        RECT  2.480 1.340 2.680 2.360 ;
        RECT  1.000 1.340 3.880 1.900 ;
        RECT  3.560 0.880 3.880 2.360 ;
        RECT  0.720 0.880 1.160 1.160 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.780 1.620 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.340 -0.280 1.980 0.640 ;
        RECT  3.040 -0.280 4.040 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.350 2.580 1.990 3.480 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVCKMHD

MACRO INVCKNHD
    CLASS CORE ;
    FOREIGN INVCKNHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.000 0.840 1.200 2.300 ;
        RECT  0.620 2.140 1.200 2.300 ;
        RECT  2.180 0.940 2.460 2.300 ;
        RECT  2.180 1.290 2.500 2.300 ;
        RECT  3.260 0.940 3.540 2.300 ;
        RECT  1.000 1.290 4.740 1.890 ;
        RECT  4.300 0.940 4.740 2.300 ;
        RECT  0.660 0.840 1.200 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.320 0.780 1.620 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.900 0.640 ;
        RECT  2.800 -0.280 5.100 0.400 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.260 2.580 1.900 3.480 ;
        RECT  2.740 2.620 3.020 3.480 ;
        RECT  3.780 2.620 4.060 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVCKNHD

MACRO INVCKQHD
    CLASS CORE ;
    FOREIGN INVCKQHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.100 0.940 9.780 2.130 ;
        RECT  0.620 1.970 9.780 2.130 ;
        RECT  0.660 0.940 9.780 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.840 1.600 ;
        RECT  0.100 1.320 0.340 1.880 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.100 -0.280 10.300 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.620 1.420 3.480 ;
        RECT  2.260 2.620 2.540 3.480 ;
        RECT  3.300 2.620 3.580 3.480 ;
        RECT  4.340 2.620 4.620 3.480 ;
        RECT  5.450 2.580 6.090 3.480 ;
        RECT  6.900 2.620 7.180 3.480 ;
        RECT  7.940 2.620 8.220 3.480 ;
        RECT  8.980 2.620 9.260 3.480 ;
        RECT  10.020 2.620 10.300 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVCKQHD

MACRO INVDHD
    CLASS CORE ;
    FOREIGN INVDHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 0.790 0.320 1.070 ;
        RECT  0.100 2.080 0.320 2.360 ;
        RECT  0.100 0.790 0.300 2.360 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        RECT  0.620 -0.280 0.900 1.010 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        RECT  0.620 2.140 0.900 3.480 ;
        END
    END VCC
END INVDHD

MACRO INVGHD
    CLASS CORE ;
    FOREIGN INVGHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 0.790 0.840 1.070 ;
        RECT  0.500 2.080 0.840 2.360 ;
        RECT  0.500 0.790 0.700 2.360 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.280 1.460 1.500 1.740 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.280 -0.280 1.440 0.820 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 0.320 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.280 2.360 1.440 3.480 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 2.360 0.320 3.480 ;
        END
    END VCC
END INVGHD

MACRO INVHHD
    CLASS CORE ;
    FOREIGN INVHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.780 1.900 2.420 ;
        RECT  0.100 2.220 1.900 2.420 ;
        RECT  0.100 0.780 1.900 0.980 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.860 -0.280 1.140 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.860 2.580 1.140 3.480 ;
        END
    END VCC
END INVHHD

MACRO INVIHD
    CLASS CORE ;
    FOREIGN INVIHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 0.900 2.300 1.180 ;
        RECT  2.080 2.020 2.300 2.300 ;
        RECT  2.100 0.900 2.300 2.300 ;
        RECT  0.980 2.100 2.300 2.300 ;
        RECT  0.980 0.900 2.300 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 -0.280 1.780 0.730 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.460 -0.280 0.740 0.730 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.480 1.780 3.480 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.460 2.480 0.740 3.480 ;
        END
    END VCC
END INVIHD

MACRO INVJHD
    CLASS CORE ;
    FOREIGN INVJHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.900 2.300 2.300 ;
        RECT  0.980 2.100 2.300 2.300 ;
        RECT  0.980 0.900 2.300 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 -0.280 1.780 0.580 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.220 -0.280 0.500 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.620 1.780 3.480 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.220 2.580 0.500 3.480 ;
        END
    END VCC
END INVJHD

MACRO INVKHD
    CLASS CORE ;
    FOREIGN INVKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.720 0.860 1.880 2.340 ;
        RECT  1.700 0.900 1.900 2.300 ;
        RECT  0.620 2.100 1.900 2.300 ;
        RECT  0.620 0.900 1.900 1.100 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  2.420 -0.280 2.700 0.780 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.620 1.420 3.480 ;
        RECT  2.420 2.420 2.700 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVKHD

MACRO INVLHD
    CLASS CORE ;
    FOREIGN INVLHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.780 2.700 2.420 ;
        RECT  0.300 2.220 2.700 2.420 ;
        RECT  0.300 0.780 2.700 0.980 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.580 ;
        RECT  3.140 -0.280 3.420 0.780 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.820 -0.280 1.100 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.620 2.140 3.480 ;
        RECT  3.140 2.420 3.420 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.820 2.620 1.100 3.480 ;
        END
    END VCC
END INVLHD

MACRO INVMHD
    CLASS CORE ;
    FOREIGN INVMHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.780 3.100 2.420 ;
        RECT  0.700 2.220 3.100 2.420 ;
        RECT  0.700 0.780 3.100 0.980 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.580 ;
        RECT  2.260 -0.280 2.540 0.580 ;
        RECT  3.540 -0.280 3.820 0.780 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.180 -0.280 0.460 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 2.620 1.500 3.480 ;
        RECT  2.260 2.620 2.540 3.480 ;
        RECT  3.540 2.420 3.820 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.180 2.620 0.460 3.480 ;
        END
    END VCC
END INVMHD

MACRO INVNHD
    CLASS CORE ;
    FOREIGN INVNHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.070 0.820 4.330 2.380 ;
        RECT  0.860 2.120 4.330 2.380 ;
        RECT  0.860 0.820 4.330 1.080 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.420 2.300 1.960 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 -0.280 1.660 0.580 ;
        RECT  2.420 -0.280 2.700 0.580 ;
        RECT  3.460 -0.280 3.740 0.580 ;
        RECT  4.740 -0.280 5.020 0.780 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.340 -0.280 0.620 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.620 1.660 3.480 ;
        RECT  2.420 2.620 2.700 3.480 ;
        RECT  3.460 2.620 3.740 3.480 ;
        RECT  4.740 2.420 5.020 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.340 2.620 0.620 3.480 ;
        END
    END VCC
END INVNHD

MACRO INVQHD
    CLASS CORE ;
    FOREIGN INVQHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.490 0.960 10.300 2.160 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.110 11.100 1.960 ;
        RECT  10.510 1.340 11.100 1.740 ;
        END
    END I
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  2.180 -0.280 2.460 0.580 ;
        RECT  3.220 -0.280 3.500 0.580 ;
        RECT  4.260 -0.280 4.540 0.580 ;
        RECT  5.300 -0.280 5.580 0.580 ;
        RECT  6.340 -0.280 6.620 0.580 ;
        RECT  7.380 -0.280 7.660 0.580 ;
        RECT  8.420 -0.280 8.700 0.580 ;
        RECT  9.460 -0.280 9.740 0.580 ;
        RECT  10.740 -0.280 11.020 0.780 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.620 1.420 3.480 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  3.220 2.620 3.500 3.480 ;
        RECT  4.260 2.620 4.540 3.480 ;
        RECT  5.300 2.620 5.580 3.480 ;
        RECT  6.340 2.620 6.620 3.480 ;
        RECT  7.380 2.620 7.660 3.480 ;
        RECT  8.420 2.620 8.700 3.480 ;
        RECT  9.460 2.620 9.740 3.480 ;
        RECT  10.740 2.420 11.020 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END INVQHD

MACRO INVTCHD
    CLASS CORE ;
    FOREIGN INVTCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.440 1.900 2.360 ;
        RECT  1.680 2.080 1.900 2.360 ;
        RECT  1.680 0.440 1.900 0.720 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.100 2.070 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.440 1.070 0.700 1.350 ;
        RECT  0.500 0.900 1.500 1.100 ;
        RECT  1.300 0.980 1.540 1.260 ;
        RECT  0.500 0.740 0.700 1.350 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.620 2.800 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.120 2.480 1.520 2.640 ;
        RECT  1.360 1.460 1.520 2.640 ;
        RECT  0.120 1.890 0.320 2.640 ;
        RECT  0.120 0.650 0.280 2.640 ;
        RECT  1.360 1.460 1.540 1.740 ;
        RECT  0.120 0.650 0.320 0.930 ;
    END
END INVTCHD

MACRO INVTEHD
    CLASS CORE ;
    FOREIGN INVTEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.440 1.900 2.360 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.920 1.460 1.080 2.680 ;
        RECT  2.500 1.460 2.700 2.680 ;
        RECT  0.920 2.520 2.700 2.680 ;
        RECT  0.890 1.460 1.080 1.740 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.120 2.300 1.400 ;
        RECT  2.100 0.780 2.300 1.400 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.820 -0.280 3.100 0.620 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.900 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.880 2.560 3.100 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.600 2.650 0.760 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.120 1.890 0.320 2.170 ;
        RECT  0.120 1.060 0.280 2.170 ;
        RECT  1.380 1.060 1.540 1.740 ;
        RECT  0.160 0.960 0.320 1.240 ;
        RECT  0.120 1.060 1.540 1.220 ;
    END
END INVTEHD

MACRO INVTHHD
    CLASS CORE ;
    FOREIGN INVTHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 0.800 5.100 2.300 ;
        RECT  4.200 2.100 5.100 2.300 ;
        RECT  4.200 0.800 5.100 1.000 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.520 2.700 2.040 ;
        RECT  2.320 1.520 2.700 1.740 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 -0.280 1.940 0.400 ;
        RECT  3.540 -0.280 3.820 0.400 ;
        RECT  4.820 -0.280 5.100 0.620 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.420 2.580 2.700 3.480 ;
        RECT  3.580 2.620 3.860 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.040 1.840 3.340 2.120 ;
        RECT  3.180 0.880 3.340 2.120 ;
        RECT  3.180 1.520 4.740 1.680 ;
        RECT  2.600 0.880 3.340 1.040 ;
        RECT  1.160 2.040 1.700 2.200 ;
        RECT  1.160 0.560 1.320 2.200 ;
        RECT  3.730 1.200 4.240 1.360 ;
        RECT  3.730 0.560 3.890 1.360 ;
        RECT  1.160 0.560 3.890 0.720 ;
        RECT  1.960 1.200 2.120 2.170 ;
        RECT  2.860 1.200 3.020 1.660 ;
        RECT  1.480 1.260 2.120 1.540 ;
        RECT  1.960 1.200 3.020 1.360 ;
        RECT  2.180 0.880 2.340 1.360 ;
        RECT  0.280 2.420 2.040 2.580 ;
        RECT  0.100 2.030 0.980 2.190 ;
        RECT  0.820 0.800 0.980 2.190 ;
        RECT  0.100 0.800 0.980 0.960 ;
    END
END INVTHHD

MACRO INVTKHD
    CLASS CORE ;
    FOREIGN INVTKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.740 5.500 2.300 ;
        RECT  4.060 2.100 5.500 2.300 ;
        RECT  4.060 0.740 5.500 0.940 ;
        END
    END O
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.520 2.700 2.040 ;
        RECT  2.320 1.520 2.700 1.740 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END E
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 -0.280 1.940 0.400 ;
        RECT  3.500 -0.280 3.780 0.400 ;
        RECT  4.580 -0.280 4.860 0.580 ;
        RECT  5.620 -0.280 5.900 0.580 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.460 2.580 2.740 3.480 ;
        RECT  3.540 2.300 3.820 3.480 ;
        RECT  4.580 2.620 4.860 3.480 ;
        RECT  5.620 2.620 5.900 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.540 2.800 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.080 1.840 3.340 2.120 ;
        RECT  3.180 0.880 3.340 2.120 ;
        RECT  3.180 1.520 4.460 1.680 ;
        RECT  2.600 0.880 3.340 1.040 ;
        RECT  1.160 2.040 1.700 2.200 ;
        RECT  1.160 0.560 1.320 2.200 ;
        RECT  3.500 1.200 4.020 1.360 ;
        RECT  3.500 0.560 3.660 1.360 ;
        RECT  1.160 0.560 3.660 0.720 ;
        RECT  1.960 1.200 2.120 2.170 ;
        RECT  2.860 1.200 3.020 1.660 ;
        RECT  1.480 1.260 2.120 1.540 ;
        RECT  1.960 1.200 3.020 1.360 ;
        RECT  2.180 0.880 2.340 1.360 ;
        RECT  1.320 2.580 2.040 2.740 ;
        RECT  0.280 2.420 1.480 2.580 ;
        RECT  0.100 2.030 0.980 2.190 ;
        RECT  0.820 0.800 0.980 2.190 ;
        RECT  0.100 0.800 0.980 0.960 ;
    END
END INVTKHD

MACRO MAO222CHD
    CLASS CORE ;
    FOREIGN MAO222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.800 3.500 2.270 ;
        RECT  3.220 2.110 3.500 2.270 ;
        RECT  3.220 0.800 3.500 0.960 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.390 1.100 1.670 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.390 1.600 1.670 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  2.430 1.390 2.630 2.260 ;
        RECT  0.100 2.060 2.630 2.260 ;
        RECT  0.100 1.220 0.300 2.260 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 -0.280 2.940 0.640 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.720 -0.280 0.880 0.680 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 2.800 2.900 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.740 2.420 3.060 2.580 ;
        RECT  2.900 0.800 3.060 2.580 ;
        RECT  2.900 1.390 3.100 1.670 ;
        RECT  1.700 0.800 3.060 0.960 ;
        RECT  0.100 0.860 1.540 1.020 ;
        RECT  0.100 0.800 0.380 1.020 ;
        RECT  0.100 2.420 1.500 2.580 ;
    END
END MAO222CHD

MACRO MAO222EHD
    CLASS CORE ;
    FOREIGN MAO222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.800 3.500 2.270 ;
        RECT  3.220 2.110 3.500 2.270 ;
        RECT  3.220 0.800 3.500 0.960 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.180 1.100 1.900 ;
        RECT  1.980 1.390 2.140 1.900 ;
        RECT  0.900 1.740 2.140 1.900 ;
        RECT  0.860 1.300 1.100 1.580 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.600 1.580 ;
        RECT  1.300 1.180 1.500 1.580 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  2.480 1.390 2.640 2.220 ;
        RECT  0.100 2.060 2.640 2.220 ;
        RECT  0.100 1.220 0.300 2.220 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 -0.280 2.940 0.580 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.740 -0.280 0.900 0.680 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.640 2.800 2.920 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.760 2.420 3.060 2.580 ;
        RECT  2.900 0.800 3.060 2.580 ;
        RECT  2.900 1.390 3.120 1.670 ;
        RECT  1.720 0.800 3.060 0.960 ;
        RECT  0.100 0.860 1.520 1.020 ;
        RECT  0.100 0.800 0.380 1.020 ;
        RECT  0.100 2.420 1.520 2.580 ;
        RECT  0.100 2.380 0.380 2.580 ;
    END
END MAO222EHD

MACRO MAO222HHD
    CLASS CORE ;
    FOREIGN MAO222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.890 2.100 4.300 2.300 ;
        RECT  3.890 0.900 4.300 1.100 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.180 1.100 1.900 ;
        RECT  1.980 1.390 2.140 1.900 ;
        RECT  0.900 1.740 2.140 1.900 ;
        RECT  0.860 1.440 1.100 1.720 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.600 1.580 ;
        RECT  1.300 1.180 1.500 1.580 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  2.480 1.390 2.640 2.220 ;
        RECT  0.100 2.060 2.640 2.220 ;
        RECT  0.100 1.220 0.300 2.220 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.600 -0.280 2.880 0.620 ;
        RECT  4.420 -0.280 4.700 0.620 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.680 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.640 2.800 2.920 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.760 2.420 3.040 2.580 ;
        RECT  2.880 0.800 3.040 2.580 ;
        RECT  2.880 1.390 3.120 1.670 ;
        RECT  1.720 0.800 3.040 0.960 ;
        RECT  0.100 0.860 1.520 1.020 ;
        RECT  0.100 0.800 0.380 1.020 ;
        RECT  0.100 2.420 1.520 2.580 ;
        RECT  0.100 2.380 0.380 2.580 ;
    END
END MAO222HHD

MACRO MAO222KHD
    CLASS CORE ;
    FOREIGN MAO222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.240 0.900 6.560 1.100 ;
        RECT  5.260 2.100 6.630 2.300 ;
        RECT  6.100 0.900 6.300 2.300 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.390 1.100 1.670 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.390 1.600 1.670 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  2.430 1.390 2.630 2.260 ;
        RECT  0.100 2.060 2.630 2.260 ;
        RECT  0.100 1.220 0.300 2.260 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.640 -0.280 2.920 0.580 ;
        RECT  3.680 -0.280 3.960 0.580 ;
        RECT  4.720 -0.280 5.000 0.580 ;
        RECT  5.760 -0.280 6.040 0.580 ;
        RECT  6.820 -0.280 7.100 0.580 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.620 2.800 2.900 3.480 ;
        RECT  3.660 2.620 3.940 3.480 ;
        RECT  4.720 2.620 5.000 3.480 ;
        RECT  5.780 2.620 6.060 3.480 ;
        RECT  6.820 2.620 7.100 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.660 2.800 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.140 2.140 5.020 2.300 ;
        RECT  4.860 0.740 5.020 2.300 ;
        RECT  4.860 1.420 5.740 1.580 ;
        RECT  4.200 0.740 5.020 0.900 ;
        RECT  3.240 2.050 3.560 2.330 ;
        RECT  3.360 0.800 3.560 2.330 ;
        RECT  3.360 1.390 3.580 1.670 ;
        RECT  3.200 0.800 3.560 1.020 ;
        RECT  1.740 2.420 3.040 2.580 ;
        RECT  2.880 0.800 3.040 2.580 ;
        RECT  2.880 1.390 3.100 1.670 ;
        RECT  1.700 0.800 3.040 0.960 ;
        RECT  0.100 0.860 1.540 1.020 ;
        RECT  0.100 0.800 0.380 1.020 ;
        RECT  0.100 2.420 1.500 2.580 ;
    END
END MAO222KHD

MACRO MAOI1CHD
    CLASS CORE ;
    FOREIGN MAOI1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 2.340 3.480 2.620 ;
        RECT  1.700 0.740 3.500 0.900 ;
        RECT  3.320 0.740 3.480 2.620 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.780 ;
        RECT  2.480 1.360 2.700 1.640 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.820 ;
        RECT  2.660 -0.280 2.940 0.580 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.100 2.620 2.380 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.160 2.320 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.540 1.980 3.140 2.140 ;
        RECT  2.980 1.360 3.140 2.140 ;
        RECT  0.540 0.680 0.700 2.140 ;
        RECT  0.540 0.680 0.940 0.840 ;
        RECT  1.540 2.300 2.940 2.460 ;
    END
END MAOI1CHD

MACRO MAOI1EHD
    CLASS CORE ;
    FOREIGN MAOI1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.680 3.900 2.460 ;
        RECT  3.680 2.180 3.900 2.460 ;
        RECT  3.680 0.680 3.900 0.960 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.660 2.360 1.940 ;
        RECT  2.100 1.600 2.300 2.140 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 -0.280 3.380 0.700 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.940 -0.280 1.220 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.330 2.620 1.610 3.480 ;
        RECT  3.160 2.520 3.320 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.160 2.240 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.520 0.860 2.680 2.360 ;
        RECT  3.360 0.860 3.520 1.640 ;
        RECT  1.940 0.860 3.520 1.020 ;
        RECT  1.770 2.520 3.000 2.680 ;
        RECT  2.840 1.360 3.000 2.680 ;
        RECT  1.770 2.300 1.930 2.680 ;
        RECT  0.540 2.300 1.930 2.460 ;
        RECT  0.540 0.660 0.700 2.460 ;
        RECT  0.100 0.660 0.700 0.820 ;
        RECT  1.420 0.540 2.840 0.700 ;
    END
END MAOI1EHD

MACRO MAOI1HHD
    CLASS CORE ;
    FOREIGN MAOI1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.500 0.760 4.300 0.960 ;
        RECT  4.100 0.760 4.300 2.300 ;
        RECT  3.440 2.100 4.300 2.300 ;
        RECT  3.500 0.740 3.780 0.960 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        RECT  1.660 1.360 1.900 1.640 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.200 2.300 1.740 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 -0.280 3.260 0.600 ;
        RECT  4.020 -0.280 4.300 0.600 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.940 -0.280 1.220 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.620 1.460 3.480 ;
        RECT  2.920 2.620 3.200 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.320 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.300 1.980 2.620 2.140 ;
        RECT  2.460 0.760 2.620 2.140 ;
        RECT  3.260 1.140 3.420 1.640 ;
        RECT  2.460 1.140 3.420 1.300 ;
        RECT  1.900 0.760 2.620 0.920 ;
        RECT  0.540 2.300 2.940 2.460 ;
        RECT  2.780 1.460 2.940 2.460 ;
        RECT  0.540 0.660 0.700 2.460 ;
        RECT  0.100 0.660 0.700 0.820 ;
        RECT  1.420 0.440 1.700 0.660 ;
        RECT  1.420 0.440 2.780 0.600 ;
    END
END MAOI1HHD

MACRO MAOI1KHD
    CLASS CORE ;
    FOREIGN MAOI1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.900 6.700 2.300 ;
        RECT  4.840 2.100 6.700 2.300 ;
        RECT  4.840 0.900 6.700 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.780 ;
        RECT  2.480 1.360 2.700 1.640 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.820 ;
        RECT  2.660 -0.280 2.940 0.580 ;
        RECT  4.320 -0.280 4.600 0.580 ;
        RECT  5.360 -0.280 5.640 0.580 ;
        RECT  6.420 -0.280 6.700 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.100 2.620 2.380 3.480 ;
        RECT  4.320 2.620 4.600 3.480 ;
        RECT  5.380 2.620 5.660 3.480 ;
        RECT  6.420 2.620 6.700 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.780 2.140 4.620 2.300 ;
        RECT  4.460 0.790 4.620 2.300 ;
        RECT  4.460 1.420 5.970 1.580 ;
        RECT  3.800 0.790 4.620 0.950 ;
        RECT  3.280 2.340 3.480 2.620 ;
        RECT  3.320 0.740 3.480 2.620 ;
        RECT  3.320 1.420 4.260 1.580 ;
        RECT  1.700 0.740 3.500 0.900 ;
        RECT  0.540 1.980 3.140 2.140 ;
        RECT  2.980 1.360 3.140 2.140 ;
        RECT  0.540 0.680 0.700 2.140 ;
        RECT  0.540 0.680 0.940 0.840 ;
        RECT  1.540 2.300 2.940 2.460 ;
    END
END MAOI1KHD

MACRO MOAI1CHD
    CLASS CORE ;
    FOREIGN MOAI1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.320 1.980 2.680 2.140 ;
        RECT  1.940 0.860 3.500 1.020 ;
        RECT  3.300 0.860 3.500 2.340 ;
        RECT  2.520 0.860 2.680 2.140 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.360 2.360 1.640 ;
        RECT  2.100 1.240 2.300 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.000 -0.280 3.280 0.600 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.940 -0.280 1.220 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.330 2.620 1.610 3.480 ;
        RECT  2.940 2.620 3.220 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.340 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.540 2.300 3.000 2.460 ;
        RECT  2.840 1.760 3.000 2.460 ;
        RECT  0.540 0.660 0.700 2.460 ;
        RECT  0.100 0.660 0.700 0.820 ;
        RECT  1.420 0.440 1.700 0.660 ;
        RECT  1.420 0.440 2.740 0.600 ;
    END
END MOAI1CHD

MACRO MOAI1EHD
    CLASS CORE ;
    FOREIGN MOAI1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.680 3.900 2.620 ;
        RECT  3.600 2.340 3.900 2.620 ;
        RECT  3.680 0.680 3.900 0.960 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.780 ;
        RECT  2.380 1.360 2.700 1.640 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.820 ;
        RECT  1.620 -0.280 1.900 0.580 ;
        RECT  3.100 -0.280 3.380 0.580 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.020 2.620 3.300 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.940 2.280 3.440 2.440 ;
        RECT  3.280 0.740 3.440 2.440 ;
        RECT  3.280 1.360 3.510 1.640 ;
        RECT  2.500 0.740 3.440 0.900 ;
        RECT  0.540 1.960 3.020 2.120 ;
        RECT  2.860 1.360 3.020 2.120 ;
        RECT  0.540 0.680 0.700 2.120 ;
        RECT  0.540 0.680 0.900 0.840 ;
        RECT  1.360 2.600 2.820 2.760 ;
        RECT  1.360 2.580 1.740 2.760 ;
    END
END MOAI1EHD

MACRO MOAI1HHD
    CLASS CORE ;
    FOREIGN MOAI1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.850 3.900 2.420 ;
        RECT  3.560 2.140 3.900 2.420 ;
        RECT  3.560 0.850 3.900 1.130 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.780 ;
        RECT  2.380 1.360 2.700 1.640 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.820 ;
        RECT  1.620 -0.280 1.900 0.580 ;
        RECT  2.980 -0.280 3.260 0.580 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.940 2.280 3.400 2.440 ;
        RECT  3.240 0.740 3.400 2.440 ;
        RECT  3.240 1.450 3.510 1.730 ;
        RECT  2.460 0.740 3.400 0.900 ;
        RECT  0.540 1.960 3.020 2.120 ;
        RECT  2.860 1.360 3.020 2.120 ;
        RECT  0.540 0.680 0.700 2.120 ;
        RECT  0.540 0.680 0.900 0.840 ;
        RECT  1.480 2.600 2.780 2.760 ;
        RECT  1.480 2.330 1.640 2.760 ;
    END
END MOAI1HHD

MACRO MOAI1KHD
    CLASS CORE ;
    FOREIGN MOAI1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.840 0.900 6.180 1.100 ;
        RECT  4.840 2.100 6.180 2.300 ;
        RECT  5.700 0.900 5.900 2.300 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.780 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.360 0.320 1.640 ;
        RECT  0.100 1.240 0.300 1.780 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.360 2.360 1.640 ;
        RECT  2.100 1.240 2.300 1.780 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 -0.280 3.260 0.600 ;
        RECT  4.320 -0.280 4.600 0.580 ;
        RECT  5.360 -0.280 5.640 0.580 ;
        RECT  6.420 -0.280 6.700 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.940 -0.280 1.220 0.820 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.330 2.620 1.610 3.480 ;
        RECT  2.940 2.620 3.220 3.480 ;
        RECT  4.320 2.620 4.600 3.480 ;
        RECT  5.380 2.620 5.660 3.480 ;
        RECT  6.420 2.620 6.700 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.100 2.340 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.540 2.140 3.820 2.360 ;
        RECT  3.640 0.790 3.800 2.360 ;
        RECT  3.640 1.420 5.340 1.580 ;
        RECT  3.460 0.790 3.800 0.950 ;
        RECT  2.320 1.980 2.680 2.140 ;
        RECT  2.520 0.860 2.680 2.140 ;
        RECT  2.520 1.320 3.480 1.480 ;
        RECT  1.940 0.860 2.680 1.020 ;
        RECT  0.540 2.300 3.000 2.460 ;
        RECT  2.840 1.760 3.000 2.460 ;
        RECT  0.540 0.660 0.700 2.460 ;
        RECT  0.100 0.660 0.700 0.820 ;
        RECT  1.420 0.440 1.700 0.660 ;
        RECT  1.420 0.440 2.740 0.600 ;
    END
END MOAI1KHD

MACRO MUX2CHD
    CLASS CORE ;
    FOREIGN MUX2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 0.710 3.500 2.440 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.300 2.700 1.800 ;
        RECT  2.460 1.390 2.700 1.670 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.700 -0.280 0.980 0.400 ;
        RECT  2.660 -0.280 2.940 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.220 2.800 3.220 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.160 2.540 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.280 3.100 2.440 ;
        RECT  2.940 1.350 3.100 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.340 2.600 1.980 2.760 ;
        RECT  1.340 2.280 1.500 2.760 ;
        RECT  0.980 2.280 1.500 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.380 1.200 ;
        RECT  1.220 0.480 1.380 1.200 ;
        RECT  1.220 0.480 2.300 0.640 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MUX2CHD

MACRO MUX2EHD
    CLASS CORE ;
    FOREIGN MUX2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.280 0.490 3.500 2.680 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.400 0.320 1.680 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.300 2.700 1.800 ;
        RECT  2.460 1.390 2.700 1.670 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 -0.280 1.320 0.400 ;
        RECT  2.510 -0.280 2.790 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.220 2.800 2.860 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.160 2.540 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.280 3.100 2.440 ;
        RECT  2.940 1.350 3.100 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.790 2.300 2.120 ;
        RECT  2.140 0.790 2.420 1.070 ;
        RECT  1.340 2.600 1.980 2.760 ;
        RECT  1.340 2.280 1.500 2.760 ;
        RECT  0.980 2.280 1.500 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.380 1.200 ;
        RECT  1.220 0.610 1.380 1.200 ;
        RECT  1.220 0.610 1.880 0.770 ;
        RECT  1.600 0.470 2.300 0.630 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MUX2EHD

MACRO MUX2HHD
    CLASS CORE ;
    FOREIGN MUX2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.740 4.700 2.460 ;
        RECT  3.900 2.260 4.700 2.460 ;
        RECT  3.900 0.740 4.700 0.940 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.210 0.700 2.430 ;
        RECT  2.080 1.300 2.240 2.430 ;
        RECT  0.500 2.270 2.240 2.430 ;
        RECT  0.480 1.340 0.700 1.620 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.120 1.680 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.150 3.500 1.670 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.380 -0.280 3.660 0.660 ;
        RECT  4.420 -0.280 4.700 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.640 -0.280 0.920 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.380 2.620 3.660 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.640 2.620 0.920 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.400 2.300 3.740 2.460 ;
        RECT  3.580 1.940 3.740 2.460 ;
        RECT  2.400 0.960 2.560 2.460 ;
        RECT  3.580 1.940 4.340 2.100 ;
        RECT  4.180 1.390 4.340 2.100 ;
        RECT  2.920 0.960 3.080 2.120 ;
        RECT  1.320 1.900 1.920 2.060 ;
        RECT  1.760 0.920 1.920 2.060 ;
        RECT  0.160 0.560 0.320 2.160 ;
        RECT  1.440 0.460 1.600 1.700 ;
        RECT  0.160 0.560 1.720 0.720 ;
        RECT  1.440 0.460 1.720 0.720 ;
    END
END MUX2HHD

MACRO MUX2KHD
    CLASS CORE ;
    FOREIGN MUX2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.740 5.900 2.460 ;
        RECT  4.060 2.260 5.900 2.460 ;
        RECT  4.060 0.740 5.900 0.940 ;
        END
    END O
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.210 0.700 2.430 ;
        RECT  2.080 1.300 2.240 2.430 ;
        RECT  0.500 2.270 2.240 2.430 ;
        RECT  0.480 1.340 0.700 1.620 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.120 1.680 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.150 3.500 1.670 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.450 -0.280 3.730 0.400 ;
        RECT  4.580 -0.280 4.860 0.580 ;
        RECT  5.620 -0.280 5.900 0.580 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  0.640 -0.280 0.920 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.460 2.800 3.740 3.480 ;
        RECT  4.580 2.620 4.860 3.480 ;
        RECT  5.620 2.620 5.900 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.640 2.620 0.920 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.400 2.300 3.900 2.460 ;
        RECT  3.740 1.940 3.900 2.460 ;
        RECT  2.400 0.960 2.560 2.460 ;
        RECT  3.740 1.940 4.680 2.100 ;
        RECT  4.520 1.390 4.680 2.100 ;
        RECT  2.920 0.960 3.080 2.120 ;
        RECT  1.320 1.900 1.920 2.060 ;
        RECT  1.760 0.920 1.920 2.060 ;
        RECT  0.160 0.560 0.320 2.160 ;
        RECT  1.440 0.460 1.600 1.700 ;
        RECT  0.160 0.560 1.720 0.720 ;
        RECT  1.440 0.460 1.720 0.720 ;
    END
END MUX2KHD

MACRO MUX3CHD
    CLASS CORE ;
    FOREIGN MUX3CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.080 0.720 6.300 2.440 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.460 1.500 1.920 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.370 3.300 1.650 ;
        RECT  2.900 1.280 3.100 1.800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.340 0.300 1.860 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.280 2.700 1.800 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.300 4.440 1.580 ;
        RECT  4.100 1.300 4.300 1.820 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.700 -0.280 0.980 0.400 ;
        RECT  2.800 -0.280 3.440 0.400 ;
        RECT  4.440 -0.280 5.740 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 2.620 2.360 3.480 ;
        RECT  3.000 2.800 3.280 3.480 ;
        RECT  5.840 2.800 6.120 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.160 2.560 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.540 1.840 4.760 2.120 ;
        RECT  4.600 0.620 4.760 2.120 ;
        RECT  5.760 0.620 5.920 1.710 ;
        RECT  4.600 0.620 5.920 0.780 ;
        RECT  3.860 2.600 5.600 2.760 ;
        RECT  5.440 1.360 5.600 2.760 ;
        RECT  5.280 1.360 5.600 1.640 ;
        RECT  1.700 2.280 5.080 2.440 ;
        RECT  4.920 0.980 5.080 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  4.920 1.900 5.280 2.180 ;
        RECT  4.920 0.980 5.340 1.140 ;
        RECT  3.780 0.440 3.940 1.720 ;
        RECT  3.780 0.440 4.140 0.600 ;
        RECT  3.460 1.880 3.840 2.100 ;
        RECT  3.460 0.880 3.620 2.100 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.180 2.600 1.800 2.760 ;
        RECT  1.180 2.130 1.340 2.760 ;
        RECT  0.980 2.130 1.340 2.290 ;
        RECT  0.980 1.040 1.140 2.290 ;
        RECT  0.980 1.040 1.380 1.200 ;
        RECT  1.220 0.480 1.380 1.200 ;
        RECT  1.220 0.480 2.300 0.640 ;
        RECT  0.620 2.450 0.900 2.610 ;
        RECT  0.620 0.720 0.780 2.610 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MUX3CHD

MACRO MUX3EHD
    CLASS CORE ;
    FOREIGN MUX3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.080 0.720 6.300 2.440 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.460 1.500 1.920 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.370 3.300 1.650 ;
        RECT  2.900 1.280 3.100 1.800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.340 0.300 1.860 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.280 2.700 1.800 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.300 4.440 1.580 ;
        RECT  4.100 1.160 4.300 1.680 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.000 -0.280 1.220 0.460 ;
        RECT  2.800 -0.280 3.080 0.400 ;
        RECT  4.440 -0.280 5.740 0.400 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 2.620 2.360 3.480 ;
        RECT  3.000 2.800 3.280 3.480 ;
        RECT  5.560 2.520 5.720 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.160 2.560 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.260 1.900 4.760 2.060 ;
        RECT  4.600 0.620 4.760 2.060 ;
        RECT  5.760 0.620 5.920 1.670 ;
        RECT  4.600 0.620 5.920 0.780 ;
        RECT  3.860 2.600 5.400 2.760 ;
        RECT  5.240 1.360 5.400 2.760 ;
        RECT  5.240 1.360 5.440 1.640 ;
        RECT  1.700 2.280 5.080 2.440 ;
        RECT  4.920 0.980 5.080 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  4.920 0.980 5.340 1.140 ;
        RECT  3.780 0.440 3.940 1.720 ;
        RECT  3.780 0.440 4.140 0.600 ;
        RECT  3.460 1.900 3.840 2.060 ;
        RECT  3.460 0.880 3.620 2.060 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.180 2.600 1.800 2.760 ;
        RECT  1.180 2.130 1.340 2.760 ;
        RECT  0.980 2.130 1.340 2.290 ;
        RECT  0.980 1.040 1.140 2.290 ;
        RECT  0.980 1.040 1.540 1.200 ;
        RECT  1.380 0.480 1.540 1.200 ;
        RECT  1.380 0.480 2.300 0.640 ;
        RECT  0.620 2.450 0.900 2.610 ;
        RECT  0.620 0.720 0.780 2.610 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MUX3EHD

MACRO MUX3HHD
    CLASS CORE ;
    FOREIGN MUX3HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 0.740 8.300 2.460 ;
        RECT  7.500 2.260 8.300 2.460 ;
        RECT  7.500 0.740 8.300 0.940 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.210 0.700 2.430 ;
        RECT  2.080 1.300 2.240 2.430 ;
        RECT  0.500 2.270 2.240 2.430 ;
        RECT  0.480 1.340 0.700 1.620 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.400 4.740 1.680 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.120 1.680 ;
        RECT  0.900 1.240 1.100 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.150 3.500 1.670 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.240 4.300 1.760 ;
        RECT  5.700 1.300 5.860 2.440 ;
        RECT  4.120 2.280 5.860 2.440 ;
        RECT  4.120 1.240 4.280 2.440 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.420 -0.280 3.700 0.400 ;
        RECT  4.260 -0.280 4.540 0.400 ;
        RECT  6.520 -0.280 7.220 0.400 ;
        RECT  8.020 -0.280 8.300 0.580 ;
        RECT  0.000 -0.280 8.400 0.280 ;
        RECT  0.640 -0.280 0.920 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.420 2.740 3.640 3.480 ;
        RECT  6.960 2.620 7.240 3.480 ;
        RECT  8.020 2.620 8.300 3.480 ;
        RECT  0.000 2.920 8.400 3.480 ;
        RECT  0.640 2.620 0.920 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.020 0.640 6.180 2.180 ;
        RECT  6.860 1.940 7.940 2.100 ;
        RECT  7.780 1.390 7.940 2.100 ;
        RECT  6.860 0.640 7.020 2.100 ;
        RECT  6.020 0.640 7.020 0.800 ;
        RECT  3.800 2.600 6.700 2.760 ;
        RECT  6.540 0.960 6.700 2.760 ;
        RECT  3.800 2.420 3.960 2.760 ;
        RECT  2.400 2.420 3.960 2.580 ;
        RECT  2.400 0.960 2.560 2.580 ;
        RECT  4.940 1.900 5.540 2.060 ;
        RECT  5.380 0.920 5.540 2.060 ;
        RECT  3.780 0.560 3.940 2.120 ;
        RECT  5.060 0.460 5.220 1.700 ;
        RECT  3.780 0.560 5.340 0.720 ;
        RECT  5.060 0.460 5.340 0.720 ;
        RECT  2.920 0.960 3.080 2.120 ;
        RECT  1.320 1.900 1.920 2.060 ;
        RECT  1.760 0.920 1.920 2.060 ;
        RECT  0.160 0.560 0.320 2.160 ;
        RECT  1.440 0.460 1.600 1.700 ;
        RECT  0.160 0.560 1.720 0.720 ;
        RECT  1.440 0.460 1.720 0.720 ;
    END
END MUX3HHD

MACRO MUX3KHD
    CLASS CORE ;
    FOREIGN MUX3KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.740 10.700 2.460 ;
        RECT  8.860 2.260 10.700 2.460 ;
        RECT  8.860 0.740 10.700 0.940 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.210 0.700 2.430 ;
        RECT  2.700 1.300 2.860 2.430 ;
        RECT  0.500 2.270 2.860 2.430 ;
        RECT  0.480 1.340 0.700 1.620 ;
        END
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.240 6.300 1.760 ;
        RECT  6.060 1.400 6.300 1.680 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.400 1.120 1.680 ;
        RECT  0.900 1.220 1.100 1.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.780 1.390 5.100 1.670 ;
        RECT  4.900 1.150 5.100 1.670 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.720 1.240 5.880 2.440 ;
        RECT  5.700 1.240 5.900 1.760 ;
        RECT  7.180 1.300 7.340 2.440 ;
        RECT  5.720 2.280 7.340 2.440 ;
        RECT  5.580 1.340 5.900 1.620 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 -0.280 1.940 0.400 ;
        RECT  3.820 -0.280 4.100 0.660 ;
        RECT  4.900 -0.280 5.180 0.400 ;
        RECT  5.740 -0.280 6.020 0.400 ;
        RECT  8.140 -0.280 8.420 0.400 ;
        RECT  9.380 -0.280 9.660 0.580 ;
        RECT  10.420 -0.280 10.700 0.580 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.540 -0.280 0.820 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 2.620 1.880 3.480 ;
        RECT  3.820 2.620 4.100 3.480 ;
        RECT  4.960 2.740 5.120 3.480 ;
        RECT  8.380 2.520 8.540 3.480 ;
        RECT  9.380 2.620 9.660 3.480 ;
        RECT  10.420 2.620 10.700 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.540 2.620 0.820 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.500 0.640 7.660 2.180 ;
        RECT  8.540 0.640 8.700 1.670 ;
        RECT  7.500 0.640 8.700 0.800 ;
        RECT  5.400 2.600 8.180 2.760 ;
        RECT  8.020 0.960 8.180 2.760 ;
        RECT  5.400 2.300 5.560 2.760 ;
        RECT  3.020 2.300 5.560 2.460 ;
        RECT  3.020 0.960 3.180 2.460 ;
        RECT  6.420 1.900 7.020 2.060 ;
        RECT  6.860 0.920 7.020 2.060 ;
        RECT  5.260 0.560 5.420 2.120 ;
        RECT  6.540 0.460 6.700 1.740 ;
        RECT  5.260 0.560 6.820 0.720 ;
        RECT  6.540 0.460 6.820 0.720 ;
        RECT  3.540 1.960 4.660 2.120 ;
        RECT  3.540 0.960 3.700 2.120 ;
        RECT  3.540 0.960 4.660 1.120 ;
        RECT  1.080 1.900 2.540 2.060 ;
        RECT  2.380 0.920 2.540 2.060 ;
        RECT  1.740 0.880 1.900 2.060 ;
        RECT  1.100 0.880 1.900 1.040 ;
        RECT  0.160 0.560 0.320 2.160 ;
        RECT  2.060 0.560 2.220 1.740 ;
        RECT  0.160 0.560 2.380 0.720 ;
        RECT  2.100 0.460 2.380 0.720 ;
    END
END MUX3KHD

MACRO MUX4CHD
    CLASS CORE ;
    FOREIGN MUX4CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.630 9.900 2.120 ;
        RECT  9.680 1.840 9.900 2.120 ;
        RECT  9.680 0.630 9.900 0.910 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.300 1.960 ;
        RECT  1.980 1.370 2.300 1.650 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.130 5.900 1.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.370 6.360 1.650 ;
        RECT  6.100 1.130 6.300 1.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.400 1.650 ;
        RECT  0.100 1.220 0.300 1.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.500 2.050 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.880 1.370 9.100 1.650 ;
        RECT  8.900 1.130 9.100 1.650 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  9.060 -0.280 9.340 0.850 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  6.540 2.800 6.820 3.480 ;
        RECT  8.620 2.800 9.320 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.100 2.360 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 2.480 9.520 2.640 ;
        RECT  9.360 1.370 9.520 2.640 ;
        RECT  7.560 0.760 7.720 2.640 ;
        RECT  7.430 0.760 7.720 0.960 ;
        RECT  8.560 0.630 8.720 2.120 ;
        RECT  8.400 1.390 8.720 1.670 ;
        RECT  8.560 0.630 8.730 0.910 ;
        RECT  8.080 0.440 8.240 2.120 ;
        RECT  4.920 1.840 5.140 2.120 ;
        RECT  4.920 0.440 5.080 2.120 ;
        RECT  8.080 0.720 8.250 1.000 ;
        RECT  5.820 0.560 6.740 0.720 ;
        RECT  6.580 0.440 8.240 0.600 ;
        RECT  4.920 0.440 5.980 0.600 ;
        RECT  3.360 2.600 6.300 2.760 ;
        RECT  6.140 2.220 6.300 2.760 ;
        RECT  3.360 0.820 3.520 2.760 ;
        RECT  6.140 2.220 7.200 2.380 ;
        RECT  7.040 0.760 7.200 2.380 ;
        RECT  3.300 0.820 3.580 0.980 ;
        RECT  6.910 0.760 7.200 0.960 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.900 5.980 2.440 ;
        RECT  4.400 0.700 4.560 2.440 ;
        RECT  5.820 1.900 6.780 2.060 ;
        RECT  6.590 0.960 6.750 2.060 ;
        RECT  6.490 0.960 6.750 1.240 ;
        RECT  5.380 1.840 5.660 2.120 ;
        RECT  5.380 0.760 5.540 2.120 ;
        RECT  5.380 0.760 5.660 0.950 ;
        RECT  0.680 0.560 0.840 2.600 ;
        RECT  3.920 0.440 4.080 2.170 ;
        RECT  0.680 0.560 2.300 0.720 ;
        RECT  2.140 0.440 4.080 0.600 ;
        RECT  1.140 2.480 2.960 2.640 ;
        RECT  2.800 0.760 2.960 2.640 ;
        RECT  1.660 0.920 1.820 2.640 ;
        RECT  1.140 0.920 1.820 1.080 ;
        RECT  2.260 2.160 2.640 2.320 ;
        RECT  2.480 0.880 2.640 2.320 ;
        RECT  2.260 0.880 2.640 1.040 ;
    END
END MUX4CHD

MACRO MUX4EHD
    CLASS CORE ;
    FOREIGN MUX4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.630 9.900 2.120 ;
        RECT  9.680 1.840 9.900 2.120 ;
        RECT  9.680 0.630 9.900 0.910 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.300 1.960 ;
        RECT  1.980 1.370 2.300 1.650 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.130 5.900 1.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.370 6.360 1.650 ;
        RECT  6.100 1.130 6.300 1.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.400 1.650 ;
        RECT  0.100 1.220 0.300 1.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.500 2.050 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.880 1.370 9.100 1.650 ;
        RECT  8.900 1.130 9.100 1.650 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  9.060 -0.280 9.340 0.860 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  6.540 2.800 6.820 3.480 ;
        RECT  8.620 2.800 9.320 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.100 2.360 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 2.480 9.520 2.640 ;
        RECT  9.360 1.370 9.520 2.640 ;
        RECT  7.560 0.780 7.720 2.640 ;
        RECT  7.430 0.780 7.720 1.000 ;
        RECT  8.560 0.640 8.720 2.120 ;
        RECT  8.400 1.390 8.720 1.670 ;
        RECT  8.560 0.640 8.730 0.920 ;
        RECT  8.080 0.440 8.240 2.120 ;
        RECT  4.920 1.840 5.140 2.120 ;
        RECT  4.920 0.440 5.080 2.120 ;
        RECT  8.080 0.720 8.250 1.000 ;
        RECT  5.820 0.560 6.740 0.720 ;
        RECT  6.580 0.440 8.240 0.600 ;
        RECT  4.920 0.440 5.980 0.600 ;
        RECT  3.370 2.600 6.300 2.760 ;
        RECT  6.140 2.220 6.300 2.760 ;
        RECT  3.370 0.820 3.530 2.760 ;
        RECT  6.140 2.220 7.200 2.380 ;
        RECT  7.040 0.780 7.200 2.380 ;
        RECT  6.910 0.780 7.200 1.000 ;
        RECT  3.300 0.820 3.580 0.980 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.900 5.980 2.440 ;
        RECT  4.400 0.700 4.560 2.440 ;
        RECT  5.820 1.900 6.780 2.060 ;
        RECT  6.590 0.960 6.750 2.060 ;
        RECT  6.490 0.960 6.750 1.240 ;
        RECT  5.380 1.840 5.660 2.120 ;
        RECT  5.380 0.760 5.540 2.120 ;
        RECT  5.380 0.760 5.660 0.970 ;
        RECT  0.680 0.560 0.840 2.600 ;
        RECT  3.920 0.440 4.080 2.170 ;
        RECT  0.680 0.560 2.300 0.720 ;
        RECT  2.140 0.440 4.080 0.600 ;
        RECT  1.140 2.480 3.000 2.640 ;
        RECT  2.840 0.760 3.000 2.640 ;
        RECT  1.660 0.920 1.820 2.640 ;
        RECT  1.140 0.920 1.820 1.080 ;
        RECT  2.800 0.760 3.000 1.040 ;
        RECT  2.260 2.160 2.640 2.320 ;
        RECT  2.480 0.880 2.640 2.320 ;
        RECT  2.260 0.880 2.640 1.040 ;
    END
END MUX4EHD

MACRO MUX4HHD
    CLASS CORE ;
    FOREIGN MUX4HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.630 9.900 2.120 ;
        RECT  9.680 1.840 9.900 2.120 ;
        RECT  9.680 0.630 9.900 0.910 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.300 1.960 ;
        RECT  1.980 1.370 2.300 1.650 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.130 5.900 1.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.370 6.360 1.650 ;
        RECT  6.100 1.130 6.300 1.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.400 1.650 ;
        RECT  0.100 1.220 0.300 1.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.500 2.050 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.880 1.370 9.100 1.650 ;
        RECT  8.900 1.130 9.100 1.650 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  9.060 -0.280 9.340 0.860 ;
        RECT  10.140 -0.280 10.420 0.860 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  6.540 2.800 6.820 3.480 ;
        RECT  8.620 2.800 9.320 3.480 ;
        RECT  10.140 2.620 10.420 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.100 2.320 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 2.480 9.520 2.640 ;
        RECT  9.360 1.370 9.520 2.640 ;
        RECT  7.560 0.780 7.720 2.640 ;
        RECT  7.430 0.780 7.720 1.000 ;
        RECT  8.560 0.640 8.720 2.120 ;
        RECT  8.400 1.390 8.720 1.670 ;
        RECT  8.560 0.640 8.730 0.920 ;
        RECT  8.080 0.440 8.240 2.120 ;
        RECT  4.920 1.840 5.140 2.120 ;
        RECT  4.920 0.440 5.080 2.120 ;
        RECT  8.080 0.720 8.250 1.000 ;
        RECT  5.820 0.560 6.740 0.720 ;
        RECT  6.580 0.440 8.240 0.600 ;
        RECT  4.920 0.440 5.980 0.600 ;
        RECT  3.370 2.600 6.300 2.760 ;
        RECT  6.140 2.220 6.300 2.760 ;
        RECT  3.370 0.820 3.530 2.760 ;
        RECT  6.140 2.220 7.200 2.380 ;
        RECT  7.040 0.780 7.200 2.380 ;
        RECT  6.910 0.780 7.200 1.000 ;
        RECT  3.300 0.820 3.580 0.980 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.900 5.980 2.440 ;
        RECT  4.400 0.700 4.560 2.440 ;
        RECT  5.820 1.900 6.780 2.060 ;
        RECT  6.590 0.960 6.750 2.060 ;
        RECT  6.490 0.960 6.750 1.240 ;
        RECT  5.380 1.840 5.660 2.120 ;
        RECT  5.380 0.760 5.540 2.120 ;
        RECT  5.380 0.760 5.660 0.970 ;
        RECT  0.680 0.560 0.840 2.560 ;
        RECT  3.920 0.440 4.080 2.170 ;
        RECT  0.680 0.560 2.300 0.720 ;
        RECT  2.140 0.440 4.080 0.600 ;
        RECT  1.140 2.480 3.000 2.640 ;
        RECT  2.840 0.760 3.000 2.640 ;
        RECT  1.660 0.920 1.820 2.640 ;
        RECT  1.140 0.920 1.820 1.080 ;
        RECT  2.800 0.760 3.000 1.040 ;
        RECT  2.260 2.160 2.640 2.320 ;
        RECT  2.480 0.880 2.640 2.320 ;
        RECT  2.260 0.880 2.640 1.040 ;
    END
END MUX4HHD

MACRO MUX4KHD
    CLASS CORE ;
    FOREIGN MUX4KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  13.700 0.900 13.900 2.300 ;
        RECT  12.040 2.100 13.900 2.300 ;
        RECT  12.040 0.900 13.900 1.100 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.300 1.960 ;
        RECT  1.980 1.370 2.300 1.650 ;
        END
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.130 5.900 1.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.370 6.360 1.650 ;
        RECT  6.100 1.130 6.300 1.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.400 1.650 ;
        RECT  0.100 1.220 0.300 1.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.500 2.050 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 1.370 10.330 1.650 ;
        RECT  10.100 1.130 10.300 1.650 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  7.580 -0.280 7.740 0.950 ;
        RECT  10.350 -0.280 10.630 0.860 ;
        RECT  11.520 -0.280 11.800 0.580 ;
        RECT  12.560 -0.280 12.840 0.580 ;
        RECT  13.620 -0.280 13.900 0.580 ;
        RECT  0.000 -0.280 14.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  6.540 2.800 6.820 3.480 ;
        RECT  7.600 2.800 7.880 3.480 ;
        RECT  9.910 2.800 10.610 3.480 ;
        RECT  11.520 2.620 11.800 3.480 ;
        RECT  12.580 2.620 12.860 3.480 ;
        RECT  13.620 2.620 13.900 3.480 ;
        RECT  0.000 2.920 14.000 3.480 ;
        RECT  0.100 2.320 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.940 2.140 11.820 2.300 ;
        RECT  11.660 0.740 11.820 2.300 ;
        RECT  11.660 1.420 13.170 1.580 ;
        RECT  11.000 0.740 11.820 0.900 ;
        RECT  8.850 2.480 10.440 2.640 ;
        RECT  10.280 1.820 10.440 2.640 ;
        RECT  8.850 0.780 9.010 2.640 ;
        RECT  10.280 1.820 11.400 1.980 ;
        RECT  11.240 1.360 11.400 1.980 ;
        RECT  8.720 0.780 9.010 0.940 ;
        RECT  9.730 1.840 10.010 2.120 ;
        RECT  9.730 0.640 9.890 2.120 ;
        RECT  9.690 1.390 9.890 1.670 ;
        RECT  9.730 0.640 10.020 0.920 ;
        RECT  9.370 0.440 9.530 2.120 ;
        RECT  7.060 1.840 7.250 2.120 ;
        RECT  7.060 0.560 7.220 2.120 ;
        RECT  7.060 1.140 8.060 1.300 ;
        RECT  7.900 0.440 8.060 1.300 ;
        RECT  9.370 0.720 9.540 1.000 ;
        RECT  7.020 0.560 7.220 0.840 ;
        RECT  7.900 0.440 9.530 0.600 ;
        RECT  8.220 0.880 8.380 2.120 ;
        RECT  3.370 2.600 6.300 2.760 ;
        RECT  6.140 2.280 6.300 2.760 ;
        RECT  3.370 0.820 3.530 2.760 ;
        RECT  6.140 2.280 7.720 2.440 ;
        RECT  7.560 1.520 7.720 2.440 ;
        RECT  7.560 1.520 8.060 1.680 ;
        RECT  3.300 0.820 3.580 0.980 ;
        RECT  4.920 1.840 5.140 2.120 ;
        RECT  4.920 0.440 5.080 2.120 ;
        RECT  5.820 0.560 6.860 0.720 ;
        RECT  6.580 0.440 6.860 0.720 ;
        RECT  4.920 0.440 5.980 0.600 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.900 5.980 2.440 ;
        RECT  4.400 0.700 4.560 2.440 ;
        RECT  5.820 1.900 6.780 2.060 ;
        RECT  6.590 0.960 6.750 2.060 ;
        RECT  6.490 0.960 6.750 1.240 ;
        RECT  5.380 1.840 5.660 2.120 ;
        RECT  5.380 0.760 5.540 2.120 ;
        RECT  5.380 0.760 5.660 0.970 ;
        RECT  0.680 0.560 0.840 2.560 ;
        RECT  3.920 0.440 4.080 2.170 ;
        RECT  0.680 0.560 2.300 0.720 ;
        RECT  2.140 0.440 4.080 0.600 ;
        RECT  1.140 2.480 3.000 2.640 ;
        RECT  2.840 0.760 3.000 2.640 ;
        RECT  1.660 0.920 1.820 2.640 ;
        RECT  1.140 2.420 1.420 2.640 ;
        RECT  1.140 0.920 1.820 1.080 ;
        RECT  2.800 0.760 3.000 1.040 ;
        RECT  2.260 2.160 2.640 2.320 ;
        RECT  2.480 0.880 2.640 2.320 ;
        RECT  2.260 0.880 2.640 1.040 ;
    END
END MUX4KHD

MACRO MUX5EHD
    CLASS CORE ;
    FOREIGN MUX5EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.900 0.630 15.100 2.120 ;
        RECT  14.780 1.840 15.100 2.120 ;
        RECT  14.780 0.630 15.100 0.910 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.300 1.960 ;
        RECT  1.980 1.370 2.300 1.650 ;
        END
    END S0
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.700 1.130 11.900 1.880 ;
        RECT  11.620 1.370 11.900 1.650 ;
        END
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.130 5.900 1.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.370 6.360 1.650 ;
        RECT  6.100 1.130 6.300 1.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.400 1.650 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END B
    PIN S2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  14.100 1.130 14.300 1.880 ;
        RECT  13.960 1.370 14.300 1.650 ;
        END
    END S2
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.320 1.500 1.880 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 1.130 10.300 1.880 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  7.530 -0.280 7.810 0.400 ;
        RECT  10.280 -0.280 10.560 0.860 ;
        RECT  11.420 -0.280 11.700 0.400 ;
        RECT  14.140 -0.280 14.420 0.900 ;
        RECT  0.000 -0.280 15.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.960 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  6.540 2.800 6.820 3.480 ;
        RECT  7.580 2.800 7.860 3.480 ;
        RECT  9.780 2.800 10.480 3.480 ;
        RECT  11.430 2.460 11.710 3.480 ;
        RECT  13.690 2.800 14.390 3.480 ;
        RECT  0.000 2.920 15.200 3.480 ;
        RECT  0.100 2.360 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  12.630 2.480 14.620 2.640 ;
        RECT  14.460 1.370 14.620 2.640 ;
        RECT  12.630 0.760 12.790 2.640 ;
        RECT  12.570 0.760 12.850 0.920 ;
        RECT  13.560 1.840 13.800 2.120 ;
        RECT  13.560 0.660 13.720 2.120 ;
        RECT  13.470 1.370 13.720 1.650 ;
        RECT  13.560 0.660 13.810 0.940 ;
        RECT  10.920 0.570 11.080 2.210 ;
        RECT  13.150 0.440 13.310 2.160 ;
        RECT  13.150 0.700 13.330 0.980 ;
        RECT  10.920 0.570 12.020 0.730 ;
        RECT  11.860 0.440 13.310 0.600 ;
        RECT  12.060 0.900 12.220 2.680 ;
        RECT  12.050 2.360 12.220 2.640 ;
        RECT  8.720 2.480 10.760 2.640 ;
        RECT  10.600 1.370 10.760 2.640 ;
        RECT  8.720 0.780 8.880 2.640 ;
        RECT  8.650 0.780 8.930 0.940 ;
        RECT  9.720 0.640 9.880 2.120 ;
        RECT  9.560 1.390 9.880 1.670 ;
        RECT  9.720 0.640 9.950 0.920 ;
        RECT  9.240 0.440 9.400 2.120 ;
        RECT  7.040 1.840 7.240 2.120 ;
        RECT  7.040 1.140 7.200 2.120 ;
        RECT  7.020 1.140 7.910 1.300 ;
        RECT  7.750 0.570 7.910 1.300 ;
        RECT  7.020 0.880 7.180 1.300 ;
        RECT  9.240 0.720 9.470 1.000 ;
        RECT  7.750 0.570 8.130 0.730 ;
        RECT  7.970 0.440 9.400 0.600 ;
        RECT  8.130 1.840 8.360 2.120 ;
        RECT  8.130 0.980 8.290 2.120 ;
        RECT  8.090 0.980 8.370 1.140 ;
        RECT  3.370 2.600 6.300 2.760 ;
        RECT  6.140 2.280 6.300 2.760 ;
        RECT  3.370 0.760 3.530 2.760 ;
        RECT  6.140 2.280 7.960 2.440 ;
        RECT  7.800 1.460 7.960 2.440 ;
        RECT  7.740 1.460 7.960 1.740 ;
        RECT  3.300 0.760 3.580 0.920 ;
        RECT  4.920 1.840 5.140 2.120 ;
        RECT  4.920 0.440 5.080 2.120 ;
        RECT  5.820 0.560 7.010 0.720 ;
        RECT  6.730 0.440 7.010 0.720 ;
        RECT  4.920 0.440 5.980 0.600 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.900 5.980 2.440 ;
        RECT  4.400 0.700 4.560 2.440 ;
        RECT  5.820 1.900 6.780 2.060 ;
        RECT  6.590 0.960 6.750 2.060 ;
        RECT  6.490 0.960 6.750 1.240 ;
        RECT  5.380 1.840 5.660 2.120 ;
        RECT  5.380 0.760 5.540 2.120 ;
        RECT  5.380 0.760 5.660 0.970 ;
        RECT  0.680 0.560 0.840 2.600 ;
        RECT  3.920 0.440 4.080 2.170 ;
        RECT  0.680 0.560 2.300 0.720 ;
        RECT  2.140 0.440 4.080 0.600 ;
        RECT  1.140 2.480 3.000 2.640 ;
        RECT  2.840 0.760 3.000 2.640 ;
        RECT  1.660 0.920 1.820 2.640 ;
        RECT  1.140 2.420 1.420 2.640 ;
        RECT  1.140 0.920 1.820 1.080 ;
        RECT  2.800 0.760 3.000 1.040 ;
        RECT  2.260 2.160 2.640 2.320 ;
        RECT  2.480 0.880 2.640 2.320 ;
        RECT  2.260 0.880 2.640 1.040 ;
    END
END MUX5EHD

MACRO MUXB2BHD
    CLASS CORE ;
    FOREIGN MUXB2BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.780 4.300 2.760 ;
        RECT  3.980 2.600 4.300 2.760 ;
        RECT  3.500 0.780 4.300 0.980 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END EB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.940 -0.280 1.220 0.400 ;
        RECT  2.860 -0.280 4.300 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.160 -0.280 0.320 0.920 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.800 2.480 3.480 ;
        RECT  3.060 2.620 3.340 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.160 2.520 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.280 3.940 2.440 ;
        RECT  3.780 1.460 3.940 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.240 2.600 1.940 2.760 ;
        RECT  1.240 2.280 1.400 2.760 ;
        RECT  0.980 2.280 1.400 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.540 1.200 ;
        RECT  1.380 0.480 1.540 1.200 ;
        RECT  1.380 0.480 2.300 0.640 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MUXB2BHD

MACRO MUXB2CHD
    CLASS CORE ;
    FOREIGN MUXB2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.810 4.300 2.760 ;
        RECT  3.980 2.600 4.300 2.760 ;
        RECT  3.500 0.810 4.300 1.010 ;
        END
    END O
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END EB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.940 -0.280 1.220 0.400 ;
        RECT  2.860 -0.280 4.300 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.160 -0.280 0.320 0.920 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.800 2.480 3.480 ;
        RECT  3.060 2.620 3.340 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.160 2.520 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.280 3.940 2.440 ;
        RECT  3.780 1.460 3.940 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.240 2.600 1.940 2.760 ;
        RECT  1.240 2.280 1.400 2.760 ;
        RECT  0.980 2.280 1.400 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.540 1.200 ;
        RECT  1.380 0.470 1.540 1.200 ;
        RECT  1.380 0.470 2.300 0.630 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MUXB2CHD

MACRO MUXB4CHD
    CLASS CORE ;
    FOREIGN MUXB4CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 1.010 10.700 1.210 ;
        RECT  10.500 1.010 10.700 2.120 ;
        RECT  10.480 1.840 10.700 2.120 ;
        RECT  9.700 0.630 9.900 1.210 ;
        END
    END O
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.370 2.300 1.960 ;
        RECT  1.980 1.370 2.300 1.650 ;
        END
    END S0
    PIN EB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 1.370 9.520 1.650 ;
        RECT  9.300 1.130 9.500 1.650 ;
        END
    END EB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.130 5.900 1.650 ;
        END
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.370 6.360 1.650 ;
        RECT  6.100 1.130 6.300 1.650 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.400 1.650 ;
        RECT  0.100 1.220 0.300 1.740 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.370 1.500 2.050 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.880 1.370 9.100 1.650 ;
        RECT  8.900 1.130 9.100 1.650 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.400 ;
        RECT  6.140 -0.280 6.420 0.400 ;
        RECT  9.060 -0.280 9.340 0.850 ;
        RECT  10.420 -0.280 10.700 0.850 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  6.540 2.800 6.820 3.480 ;
        RECT  9.080 2.800 9.360 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.100 2.360 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.560 2.480 10.280 2.640 ;
        RECT  10.120 1.460 10.280 2.640 ;
        RECT  7.560 0.780 7.720 2.640 ;
        RECT  7.430 0.780 7.720 1.000 ;
        RECT  8.560 0.630 8.720 2.160 ;
        RECT  8.400 1.390 8.720 1.670 ;
        RECT  8.560 0.630 8.730 0.910 ;
        RECT  8.080 0.440 8.240 2.120 ;
        RECT  4.920 1.840 5.140 2.120 ;
        RECT  4.920 0.440 5.080 2.120 ;
        RECT  8.080 0.720 8.250 1.000 ;
        RECT  5.820 0.560 6.740 0.720 ;
        RECT  6.580 0.440 8.240 0.600 ;
        RECT  4.920 0.440 5.980 0.600 ;
        RECT  3.380 2.600 6.300 2.760 ;
        RECT  6.140 2.220 6.300 2.760 ;
        RECT  3.380 0.820 3.540 2.760 ;
        RECT  6.140 2.220 7.200 2.380 ;
        RECT  7.040 0.780 7.200 2.380 ;
        RECT  6.910 0.780 7.200 1.000 ;
        RECT  3.300 0.820 3.580 0.980 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.900 5.980 2.440 ;
        RECT  4.400 0.700 4.560 2.440 ;
        RECT  5.820 1.900 6.780 2.060 ;
        RECT  6.590 0.960 6.750 2.060 ;
        RECT  6.490 0.960 6.750 1.240 ;
        RECT  5.380 1.840 5.660 2.120 ;
        RECT  5.380 0.760 5.540 2.120 ;
        RECT  5.380 0.760 5.660 0.970 ;
        RECT  0.680 0.560 0.840 2.600 ;
        RECT  3.920 0.440 4.080 2.170 ;
        RECT  0.680 0.560 2.300 0.720 ;
        RECT  2.140 0.440 4.080 0.600 ;
        RECT  1.140 2.480 2.960 2.640 ;
        RECT  2.800 0.760 2.960 2.640 ;
        RECT  2.800 2.240 3.000 2.520 ;
        RECT  1.660 0.920 1.820 2.640 ;
        RECT  1.140 0.920 1.820 1.080 ;
        RECT  2.260 2.160 2.640 2.320 ;
        RECT  2.480 0.900 2.640 2.320 ;
        RECT  2.260 0.900 2.640 1.060 ;
    END
END MUXB4CHD

MACRO MXL2CHD
    CLASS CORE ;
    FOREIGN MXL2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.600 3.500 2.380 ;
        RECT  2.700 2.220 3.500 2.380 ;
        RECT  2.140 0.600 3.500 0.760 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.220 1.100 1.740 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.740 ;
        RECT  1.620 1.340 1.900 1.620 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.220 2.700 1.740 ;
        RECT  2.420 1.340 2.700 1.620 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.220 -0.280 3.500 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.620 1.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.180 2.600 3.500 2.760 ;
        RECT  3.220 2.540 3.500 2.760 ;
        RECT  1.240 2.300 1.400 2.650 ;
        RECT  2.180 2.300 2.340 2.760 ;
        RECT  1.240 2.300 2.340 2.460 ;
        RECT  0.160 0.880 0.320 2.160 ;
        RECT  0.160 1.900 3.140 2.060 ;
        RECT  2.980 1.370 3.140 2.060 ;
    END
END MXL2CHD

MACRO MXL2EHD
    CLASS CORE ;
    FOREIGN MXL2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 0.600 4.700 2.680 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.390 2.760 1.670 ;
        RECT  2.500 1.240 2.700 1.740 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.700 -0.280 0.980 0.400 ;
        RECT  2.660 -0.280 2.940 0.400 ;
        RECT  3.920 -0.280 4.080 1.180 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.220 2.800 2.860 3.480 ;
        RECT  3.920 2.020 4.080 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.160 2.540 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.440 0.840 3.600 2.320 ;
        RECT  3.440 1.400 4.310 1.560 ;
        RECT  1.700 2.280 3.260 2.440 ;
        RECT  3.100 1.390 3.260 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.140 1.900 2.460 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.340 2.600 1.980 2.760 ;
        RECT  1.340 2.280 1.500 2.760 ;
        RECT  0.980 2.280 1.500 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.380 1.200 ;
        RECT  1.220 0.480 1.380 1.200 ;
        RECT  1.220 0.480 2.300 0.640 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MXL2EHD

MACRO MXL2HHD
    CLASS CORE ;
    FOREIGN MXL2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.740 5.500 2.360 ;
        RECT  4.700 2.160 5.500 2.360 ;
        RECT  4.700 0.740 5.500 0.940 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.940 -0.280 1.220 0.400 ;
        RECT  3.090 -0.280 3.370 0.400 ;
        RECT  4.200 -0.280 4.360 1.180 ;
        RECT  5.220 -0.280 5.500 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.800 2.480 3.480 ;
        RECT  3.100 2.800 3.380 3.480 ;
        RECT  4.200 2.020 4.360 3.480 ;
        RECT  5.220 2.620 5.500 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.160 2.430 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.720 0.710 3.880 2.460 ;
        RECT  3.720 1.400 4.590 1.560 ;
        RECT  1.700 2.280 3.540 2.440 ;
        RECT  3.380 1.390 3.540 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.140 1.900 2.460 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.240 2.600 1.940 2.760 ;
        RECT  1.240 2.280 1.400 2.760 ;
        RECT  0.980 2.280 1.400 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.540 1.200 ;
        RECT  1.380 0.480 1.540 1.200 ;
        RECT  1.380 0.480 2.300 0.640 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MXL2HHD

MACRO MXL2KHD
    CLASS CORE ;
    FOREIGN MXL2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 0.740 6.700 2.360 ;
        RECT  4.860 2.160 6.700 2.360 ;
        RECT  4.860 0.740 6.700 0.940 ;
        END
    END OB
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.400 1.540 1.680 ;
        RECT  1.300 1.400 1.500 1.920 ;
        END
    END S
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.760 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.940 -0.280 1.220 0.400 ;
        RECT  3.090 -0.280 3.370 0.400 ;
        RECT  4.360 -0.280 4.520 1.220 ;
        RECT  5.380 -0.280 5.660 0.580 ;
        RECT  6.420 -0.280 6.700 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.800 2.480 3.480 ;
        RECT  3.100 2.800 3.380 3.480 ;
        RECT  4.360 2.020 4.520 3.480 ;
        RECT  5.380 2.620 5.660 3.480 ;
        RECT  6.420 2.620 6.700 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.160 2.540 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.720 0.920 3.880 2.300 ;
        RECT  3.720 1.400 4.750 1.560 ;
        RECT  1.700 2.280 3.540 2.440 ;
        RECT  3.380 1.390 3.540 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  2.260 0.800 2.420 2.120 ;
        RECT  1.240 2.600 1.940 2.760 ;
        RECT  1.240 2.280 1.400 2.760 ;
        RECT  0.980 2.280 1.400 2.440 ;
        RECT  0.980 1.040 1.140 2.440 ;
        RECT  0.980 1.040 1.540 1.200 ;
        RECT  1.380 0.460 1.540 1.200 ;
        RECT  1.380 0.460 2.300 0.620 ;
        RECT  0.620 2.600 0.900 2.760 ;
        RECT  0.620 0.720 0.780 2.760 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MXL2KHD

MACRO MXL3EHD
    CLASS CORE ;
    FOREIGN MXL3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.460 1.500 1.920 ;
        END
    END S0
    PIN OB
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.880 0.600 7.100 2.730 ;
        END
    END OB
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.370 3.300 1.650 ;
        RECT  2.900 1.280 3.100 1.800 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.340 0.300 1.860 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.280 2.700 1.800 ;
        END
    END A
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 1.300 4.440 1.580 ;
        RECT  4.100 1.300 4.300 1.820 ;
        END
    END S1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.700 -0.280 0.980 0.400 ;
        RECT  2.800 -0.280 3.440 0.400 ;
        RECT  4.440 -0.280 6.540 0.400 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.160 -0.280 0.320 0.940 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 2.620 2.360 3.480 ;
        RECT  3.000 2.800 3.280 3.480 ;
        RECT  5.790 2.800 6.430 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.160 2.560 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.760 2.280 6.720 2.440 ;
        RECT  6.560 1.390 6.720 2.440 ;
        RECT  5.760 0.960 5.920 2.440 ;
        RECT  4.540 1.840 4.760 2.120 ;
        RECT  4.600 0.620 4.760 2.120 ;
        RECT  6.080 0.620 6.240 1.670 ;
        RECT  4.600 0.620 6.240 0.780 ;
        RECT  3.860 2.600 5.600 2.760 ;
        RECT  5.440 1.360 5.600 2.760 ;
        RECT  5.280 1.360 5.600 1.640 ;
        RECT  1.700 2.280 5.120 2.440 ;
        RECT  4.960 0.980 5.120 2.440 ;
        RECT  1.700 0.960 1.860 2.440 ;
        RECT  4.960 1.900 5.280 2.180 ;
        RECT  4.960 0.980 5.340 1.140 ;
        RECT  3.780 0.440 3.940 1.720 ;
        RECT  3.780 0.440 4.140 0.600 ;
        RECT  3.460 1.900 3.880 2.060 ;
        RECT  3.460 0.880 3.620 2.060 ;
        RECT  2.140 1.960 2.500 2.120 ;
        RECT  2.140 0.800 2.300 2.120 ;
        RECT  2.140 0.800 2.420 1.080 ;
        RECT  1.180 2.600 1.800 2.760 ;
        RECT  1.180 2.130 1.340 2.760 ;
        RECT  0.980 2.130 1.340 2.290 ;
        RECT  0.980 1.040 1.140 2.290 ;
        RECT  0.980 1.040 1.380 1.200 ;
        RECT  1.220 0.480 1.380 1.200 ;
        RECT  1.220 0.480 2.300 0.640 ;
        RECT  0.620 2.450 0.900 2.610 ;
        RECT  0.620 0.720 0.780 2.610 ;
        RECT  0.620 0.720 0.900 0.880 ;
    END
END MXL3EHD

MACRO ND2CHD
    CLASS CORE ;
    FOREIGN ND2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 0.700 0.700 2.360 ;
        RECT  0.500 2.080 0.840 2.360 ;
        RECT  0.100 0.700 0.700 0.900 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.900 1.500 1.960 ;
        RECT  1.280 1.340 1.500 1.620 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.110 0.300 1.960 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  1.140 -0.280 1.420 0.680 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.220 1.420 3.480 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 2.160 0.340 3.480 ;
        END
    END VCC
END ND2CHD

MACRO ND2DHD
    CLASS CORE ;
    FOREIGN ND2DHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 0.700 0.700 2.360 ;
        RECT  0.500 2.080 0.840 2.360 ;
        RECT  0.100 0.700 0.700 0.900 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.900 1.500 1.960 ;
        RECT  1.280 1.340 1.500 1.620 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.110 0.300 1.960 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  1.140 -0.280 1.420 0.740 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.320 1.420 3.480 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 2.320 0.340 3.480 ;
        END
    END VCC
END ND2DHD

MACRO ND2HHD
    CLASS CORE ;
    FOREIGN ND2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.620 2.160 0.900 2.320 ;
        RECT  0.620 2.520 0.900 2.680 ;
        RECT  1.720 2.000 1.880 2.660 ;
        RECT  1.680 0.920 2.700 1.080 ;
        RECT  0.680 2.120 2.700 2.280 ;
        RECT  2.500 0.920 2.700 2.280 ;
        RECT  0.680 2.120 0.840 2.680 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.240 1.240 1.960 1.590 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.640 -0.280 0.920 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.560 1.420 3.480 ;
        RECT  2.180 2.440 2.460 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.200 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.080 0.800 1.380 0.960 ;
        RECT  1.220 0.600 1.380 0.960 ;
        RECT  1.220 0.600 2.480 0.760 ;
    END
END ND2HHD

MACRO ND2KHD
    CLASS CORE ;
    FOREIGN ND2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 2.060 1.420 2.220 ;
        RECT  0.940 0.460 1.220 1.000 ;
        RECT  1.140 2.060 1.420 2.680 ;
        RECT  2.180 2.100 2.460 2.680 ;
        RECT  2.820 0.460 3.100 1.000 ;
        RECT  3.220 2.100 3.500 2.680 ;
        RECT  1.140 2.100 4.700 2.300 ;
        RECT  0.940 0.800 4.700 1.000 ;
        RECT  4.400 0.800 4.700 2.660 ;
        RECT  4.260 2.020 4.700 2.660 ;
        RECT  0.100 2.060 0.380 2.450 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.140 0.320 1.420 ;
        RECT  3.540 1.460 3.700 1.880 ;
        RECT  0.100 1.720 3.700 1.880 ;
        RECT  0.100 0.840 0.300 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.760 1.180 3.280 1.500 ;
        RECT  1.700 1.180 1.900 1.560 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.880 -0.280 2.160 0.580 ;
        RECT  3.660 -0.280 3.940 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.660 2.540 1.940 3.480 ;
        RECT  2.700 2.540 2.980 3.480 ;
        RECT  3.740 2.540 4.020 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.620 2.380 0.900 3.480 ;
        END
    END VCC
END ND2KHD

MACRO ND3CHD
    CLASS CORE ;
    FOREIGN ND3CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.740 2.120 2.020 2.340 ;
        RECT  1.460 0.500 2.300 0.700 ;
        RECT  2.100 0.500 2.300 2.320 ;
        RECT  0.620 2.120 2.300 2.320 ;
        RECT  1.460 0.500 1.740 0.860 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 1.460 1.100 1.740 ;
        RECT  0.900 1.220 1.100 1.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.220 1.900 1.960 ;
        RECT  1.380 1.460 1.900 1.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.540 1.740 ;
        RECT  0.100 1.220 0.300 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.140 -0.280 0.420 0.870 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.480 1.460 3.480 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.100 2.260 0.380 3.480 ;
        END
    END VCC
END ND3CHD

MACRO ND3EHD
    CLASS CORE ;
    FOREIGN ND3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.660 1.980 1.940 2.280 ;
        RECT  1.460 0.480 2.700 0.680 ;
        RECT  2.500 0.480 2.700 1.140 ;
        RECT  2.700 1.980 2.980 2.280 ;
        RECT  2.500 0.940 3.500 1.140 ;
        RECT  3.300 0.940 3.500 2.140 ;
        RECT  0.620 1.980 3.500 2.140 ;
        RECT  0.620 1.980 0.900 2.280 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.780 1.340 1.100 1.500 ;
        RECT  0.900 0.840 1.100 1.500 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.590 1.300 1.940 1.500 ;
        RECT  1.700 0.840 1.900 1.500 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.820 ;
        RECT  2.840 1.520 3.120 1.820 ;
        RECT  0.100 1.660 3.120 1.820 ;
        RECT  0.100 0.840 0.300 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.140 -0.280 3.420 0.780 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.300 1.420 3.480 ;
        RECT  2.180 2.300 2.460 3.480 ;
        RECT  3.220 2.300 3.500 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.300 0.380 3.480 ;
        END
    END VCC
END ND3EHD

MACRO ND3HHD
    CLASS CORE ;
    FOREIGN ND3HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.540 2.100 3.740 2.740 ;
        RECT  3.540 0.900 4.300 1.100 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.540 2.100 4.300 2.300 ;
        RECT  3.540 0.440 3.740 1.100 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 1.460 1.100 1.740 ;
        RECT  0.900 0.840 1.100 1.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.380 1.460 1.900 1.740 ;
        RECT  1.700 0.840 1.900 1.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.540 1.740 ;
        RECT  0.100 1.220 0.300 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 -0.280 3.260 0.860 ;
        RECT  4.020 -0.280 4.300 0.720 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.140 -0.280 0.420 0.730 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.320 1.420 3.480 ;
        RECT  2.980 2.240 3.260 3.480 ;
        RECT  4.020 2.510 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.250 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.520 0.780 2.680 2.640 ;
        RECT  2.520 1.440 3.700 1.600 ;
        RECT  1.700 1.940 1.900 2.420 ;
        RECT  0.660 1.940 0.860 2.420 ;
        RECT  0.660 1.940 2.300 2.140 ;
        RECT  2.100 0.440 2.300 2.140 ;
        RECT  1.460 0.440 2.300 0.640 ;
    END
END ND3HHD

MACRO ND4CHD
    CLASS CORE ;
    FOREIGN ND4CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.420 1.980 4.700 2.260 ;
        RECT  4.500 0.840 4.700 2.360 ;
        RECT  4.420 0.840 4.700 1.120 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.180 1.540 1.460 ;
        RECT  1.300 1.100 1.500 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.180 2.300 1.960 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.100 1.960 ;
        RECT  0.880 1.340 1.100 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.740 0.320 2.020 ;
        RECT  0.100 1.240 0.300 2.030 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.280 2.600 0.700 ;
        RECT  3.360 -0.280 3.640 0.760 ;
        RECT  3.840 -0.280 4.120 1.040 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.940 -0.280 1.220 0.880 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.660 1.460 3.480 ;
        RECT  2.320 2.660 2.600 3.480 ;
        RECT  3.840 2.060 4.120 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.220 0.360 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.420 0.920 3.580 2.650 ;
        RECT  3.420 1.460 4.080 1.620 ;
        RECT  3.040 0.920 3.580 1.080 ;
        RECT  3.040 0.540 3.200 1.080 ;
        RECT  2.840 0.540 3.200 0.700 ;
        RECT  1.740 0.860 1.900 2.180 ;
        RECT  2.720 1.400 3.260 1.560 ;
        RECT  2.720 0.860 2.880 1.560 ;
        RECT  1.740 0.860 2.880 1.020 ;
        RECT  1.900 0.480 2.060 1.020 ;
        RECT  0.520 2.340 2.880 2.500 ;
        RECT  2.720 1.820 2.880 2.500 ;
        RECT  0.520 2.280 0.900 2.500 ;
        RECT  0.520 0.720 0.680 2.500 ;
        RECT  0.100 0.720 0.680 0.880 ;
    END
END ND4CHD

MACRO ND4EHD
    CLASS CORE ;
    FOREIGN ND4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.420 1.980 4.700 2.620 ;
        RECT  4.500 0.480 4.700 2.760 ;
        RECT  4.420 0.480 4.700 1.120 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.180 1.540 1.460 ;
        RECT  1.300 1.100 1.500 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.180 2.300 1.960 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.100 1.960 ;
        RECT  0.880 1.340 1.100 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.740 0.320 2.020 ;
        RECT  0.100 1.240 0.300 2.030 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.280 2.600 0.700 ;
        RECT  3.360 -0.280 3.640 0.760 ;
        RECT  3.840 -0.280 4.120 0.940 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.940 -0.280 1.220 0.880 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.640 1.460 3.480 ;
        RECT  2.320 2.640 2.600 3.480 ;
        RECT  3.840 2.260 4.120 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.220 0.360 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.420 2.370 3.620 2.650 ;
        RECT  3.460 0.920 3.620 2.650 ;
        RECT  3.460 1.460 4.080 1.620 ;
        RECT  3.040 0.920 3.620 1.080 ;
        RECT  3.040 0.540 3.200 1.080 ;
        RECT  2.840 0.540 3.200 0.700 ;
        RECT  1.740 0.860 1.900 2.160 ;
        RECT  2.720 1.320 3.300 1.480 ;
        RECT  2.720 0.860 2.880 1.480 ;
        RECT  1.740 0.860 2.880 1.020 ;
        RECT  1.900 0.480 2.060 1.020 ;
        RECT  0.520 2.320 2.880 2.480 ;
        RECT  2.720 1.740 2.880 2.480 ;
        RECT  0.520 2.280 0.900 2.480 ;
        RECT  0.520 0.720 0.680 2.480 ;
        RECT  0.100 0.720 0.680 0.880 ;
    END
END ND4EHD

MACRO ND4HHD
    CLASS CORE ;
    FOREIGN ND4HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.480 4.700 2.620 ;
        RECT  4.420 1.980 4.700 2.620 ;
        RECT  4.320 0.480 4.700 1.120 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.200 1.540 1.480 ;
        RECT  1.300 1.100 1.500 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.180 2.300 1.960 ;
        RECT  2.080 1.270 2.300 1.550 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.100 1.960 ;
        RECT  0.880 1.340 1.100 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.740 0.320 2.020 ;
        RECT  0.100 1.240 0.300 2.030 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.280 2.600 0.700 ;
        RECT  3.740 -0.280 4.020 0.940 ;
        RECT  5.060 -0.280 5.340 0.880 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.940 -0.280 1.220 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.650 1.460 3.480 ;
        RECT  2.280 2.650 2.560 3.480 ;
        RECT  3.840 2.090 4.120 3.480 ;
        RECT  5.140 2.120 5.420 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.100 2.220 0.360 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.420 0.540 3.580 2.620 ;
        RECT  3.420 1.460 4.080 1.620 ;
        RECT  2.840 0.540 3.580 0.700 ;
        RECT  1.740 0.860 1.900 2.160 ;
        RECT  2.720 1.100 3.260 1.260 ;
        RECT  2.720 0.860 2.880 1.260 ;
        RECT  1.740 0.860 2.880 1.020 ;
        RECT  1.900 0.460 2.060 1.020 ;
        RECT  0.520 2.330 2.720 2.490 ;
        RECT  2.560 1.460 2.720 2.490 ;
        RECT  0.520 2.280 0.900 2.490 ;
        RECT  0.520 0.790 0.680 2.490 ;
        RECT  0.100 0.790 0.680 0.950 ;
    END
END ND4HHD

MACRO ND4KHD
    CLASS CORE ;
    FOREIGN ND4KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.750 1.780 5.030 2.620 ;
        RECT  4.990 0.480 5.190 2.040 ;
        RECT  4.990 1.700 6.300 1.900 ;
        RECT  5.990 0.480 6.300 1.120 ;
        RECT  6.100 0.480 6.300 2.760 ;
        RECT  5.760 1.700 6.300 2.760 ;
        RECT  4.980 0.480 5.190 1.120 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.280 1.540 1.560 ;
        RECT  1.300 1.100 1.500 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.180 2.300 1.960 ;
        RECT  2.080 1.270 2.300 1.550 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.100 1.960 ;
        RECT  0.880 1.340 1.100 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.640 0.320 1.920 ;
        RECT  0.100 1.240 0.300 2.030 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.280 2.600 0.580 ;
        RECT  3.360 -0.280 3.640 0.580 ;
        RECT  4.400 -0.280 4.680 0.580 ;
        RECT  5.450 -0.280 5.730 1.120 ;
        RECT  6.570 -0.280 6.790 1.000 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.940 -0.280 1.220 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.180 2.680 1.460 3.480 ;
        RECT  2.280 2.680 2.560 3.480 ;
        RECT  4.090 2.090 4.370 3.480 ;
        RECT  5.220 2.260 5.500 3.480 ;
        RECT  6.540 2.180 6.820 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.100 2.320 0.360 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.160 1.900 3.520 2.060 ;
        RECT  3.360 0.820 3.520 2.060 ;
        RECT  4.470 1.460 4.830 1.620 ;
        RECT  4.470 0.820 4.630 1.620 ;
        RECT  2.840 0.820 4.630 0.980 ;
        RECT  3.940 0.530 4.100 0.980 ;
        RECT  2.840 0.480 3.120 0.980 ;
        RECT  0.520 2.330 2.720 2.490 ;
        RECT  2.560 1.460 2.720 2.490 ;
        RECT  3.720 1.520 3.880 2.440 ;
        RECT  2.560 2.280 3.880 2.440 ;
        RECT  0.520 2.280 0.900 2.490 ;
        RECT  0.520 0.790 0.680 2.490 ;
        RECT  3.720 1.520 4.210 1.680 ;
        RECT  0.100 0.790 0.680 0.950 ;
        RECT  1.740 0.760 1.900 2.160 ;
        RECT  3.040 1.140 3.200 1.680 ;
        RECT  2.460 1.140 3.200 1.300 ;
        RECT  2.460 0.760 2.620 1.300 ;
        RECT  1.740 0.760 2.620 0.920 ;
        RECT  1.900 0.460 2.060 0.920 ;
    END
END ND4KHD

MACRO ND5EHD
    CLASS CORE ;
    FOREIGN ND5EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.440 5.500 2.760 ;
        RECT  5.040 1.840 5.500 2.760 ;
        RECT  5.040 0.440 5.500 1.080 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.820 1.460 1.100 1.740 ;
        RECT  0.900 1.240 1.100 1.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.340 1.740 ;
        RECT  0.100 1.240 0.300 1.740 ;
        END
    END I1
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.060 1.620 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.220 3.100 1.960 ;
        RECT  2.780 1.340 3.100 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.760 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.060 -0.280 3.340 0.700 ;
        RECT  4.520 -0.280 4.740 1.000 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  1.460 -0.280 1.740 0.660 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.540 1.980 3.480 ;
        RECT  2.980 2.540 3.260 3.480 ;
        RECT  4.520 2.200 4.740 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.620 2.320 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.040 2.080 4.340 2.720 ;
        RECT  4.180 0.890 4.340 2.720 ;
        RECT  4.180 1.340 4.500 1.620 ;
        RECT  3.680 0.890 4.340 1.050 ;
        RECT  3.680 0.730 3.840 1.050 ;
        RECT  1.200 1.960 1.360 2.440 ;
        RECT  0.160 1.960 0.320 2.440 ;
        RECT  1.200 2.220 3.860 2.380 ;
        RECT  3.700 1.460 3.860 2.380 ;
        RECT  0.160 1.960 1.360 2.120 ;
        RECT  0.500 0.660 0.660 2.120 ;
        RECT  3.860 1.340 4.020 1.620 ;
        RECT  0.160 0.660 0.660 0.820 ;
        RECT  0.160 0.540 0.320 0.820 ;
        RECT  2.270 1.900 2.550 2.060 ;
        RECT  2.330 0.900 2.490 2.060 ;
        RECT  3.350 1.460 3.540 1.780 ;
        RECT  3.360 0.900 3.520 1.780 ;
        RECT  2.330 0.900 3.520 1.060 ;
    END
END ND5EHD

MACRO ND5HHD
    CLASS CORE ;
    FOREIGN ND5HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.660 5.500 2.760 ;
        RECT  5.040 1.970 5.500 2.760 ;
        RECT  5.040 0.660 5.500 0.940 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.840 1.460 1.100 1.740 ;
        RECT  0.900 0.840 1.100 1.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.340 1.740 ;
        RECT  0.100 0.840 0.300 1.740 ;
        END
    END I1
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.060 1.620 ;
        RECT  1.700 1.240 1.900 1.960 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.220 3.100 1.960 ;
        RECT  2.780 1.340 3.100 1.620 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.840 1.500 1.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.060 -0.280 3.340 0.700 ;
        RECT  4.520 -0.280 4.740 1.000 ;
        RECT  5.680 -0.280 5.900 1.000 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  1.460 -0.280 1.740 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.540 1.980 3.480 ;
        RECT  2.980 2.540 3.260 3.480 ;
        RECT  4.520 2.200 4.740 3.480 ;
        RECT  5.660 2.200 5.880 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.620 2.320 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.040 2.080 4.340 2.720 ;
        RECT  4.180 0.960 4.340 2.720 ;
        RECT  4.180 1.340 4.780 1.620 ;
        RECT  3.750 0.960 4.340 1.120 ;
        RECT  3.750 0.600 4.030 1.120 ;
        RECT  1.200 2.000 1.360 2.440 ;
        RECT  0.160 2.000 0.320 2.440 ;
        RECT  1.200 2.220 3.860 2.380 ;
        RECT  3.700 1.460 3.860 2.380 ;
        RECT  0.160 2.000 1.360 2.160 ;
        RECT  0.500 0.520 0.660 2.160 ;
        RECT  3.860 1.340 4.020 1.620 ;
        RECT  0.080 0.520 0.660 0.680 ;
        RECT  2.270 1.900 2.550 2.060 ;
        RECT  2.330 0.900 2.490 2.060 ;
        RECT  3.350 1.460 3.540 1.780 ;
        RECT  3.360 0.900 3.520 1.780 ;
        RECT  2.330 0.900 3.520 1.060 ;
    END
END ND5HHD

MACRO ND6EHD
    CLASS CORE ;
    FOREIGN ND6EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.660 5.900 2.760 ;
        RECT  5.620 2.000 5.900 2.760 ;
        RECT  5.440 0.660 5.900 0.940 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.840 ;
        RECT  0.820 1.460 1.100 1.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.340 1.740 ;
        RECT  0.100 1.240 0.300 1.740 ;
        END
    END I1
    PIN I6
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.060 1.620 ;
        RECT  1.700 1.240 1.900 1.840 ;
        END
    END I6
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.450 1.660 2.730 1.820 ;
        RECT  2.500 1.240 2.700 1.820 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.460 3.360 1.740 ;
        RECT  2.900 1.240 3.100 1.740 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.840 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.460 -0.280 3.740 0.700 ;
        RECT  4.770 -0.280 5.050 0.640 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  1.460 -0.280 1.740 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.680 1.980 3.480 ;
        RECT  2.830 2.680 3.110 3.480 ;
        RECT  3.740 2.620 4.020 3.480 ;
        RECT  5.160 2.200 5.380 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.620 2.320 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.680 1.860 4.840 2.720 ;
        RECT  4.680 1.860 5.140 2.020 ;
        RECT  4.980 0.980 5.140 2.020 ;
        RECT  4.080 0.910 4.240 1.190 ;
        RECT  4.080 0.980 5.140 1.140 ;
        RECT  1.200 2.360 3.040 2.520 ;
        RECT  4.260 1.460 4.420 2.460 ;
        RECT  0.160 2.000 0.320 2.440 ;
        RECT  2.880 2.300 4.420 2.460 ;
        RECT  1.200 2.000 1.360 2.520 ;
        RECT  0.160 2.000 1.360 2.160 ;
        RECT  0.500 0.660 0.660 2.160 ;
        RECT  4.260 1.460 4.660 1.620 ;
        RECT  4.500 1.340 4.660 1.620 ;
        RECT  0.100 0.660 0.660 0.820 ;
        RECT  2.270 1.980 2.550 2.200 ;
        RECT  2.270 1.980 3.920 2.140 ;
        RECT  3.760 0.860 3.920 2.140 ;
        RECT  3.040 0.860 3.920 1.020 ;
        RECT  3.040 0.620 3.200 1.020 ;
    END
END ND6EHD

MACRO ND8DHD
    CLASS CORE ;
    FOREIGN ND8DHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.260 0.460 8.460 1.100 ;
        RECT  8.260 0.900 8.700 1.100 ;
        RECT  8.500 0.900 8.700 2.300 ;
        RECT  7.940 2.050 8.700 2.300 ;
        RECT  7.940 2.050 8.140 2.690 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.880 ;
        RECT  1.420 1.340 1.900 1.620 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.960 ;
        END
    END I1
    PIN I8
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.940 1.620 ;
        RECT  3.700 1.240 3.900 1.960 ;
        END
    END I8
    PIN I7
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.240 4.700 1.960 ;
        END
    END I7
    PIN I6
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.240 6.300 1.960 ;
        RECT  5.980 1.340 6.300 1.620 ;
        END
    END I6
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.340 5.140 1.620 ;
        RECT  4.900 1.240 5.100 1.960 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.960 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.340 2.760 1.620 ;
        RECT  2.500 1.240 2.700 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.620 ;
        RECT  3.470 -0.280 3.750 0.780 ;
        RECT  5.760 -0.280 6.040 0.620 ;
        RECT  7.290 -0.280 7.570 0.940 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.720 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.140 2.680 2.420 3.480 ;
        RECT  3.540 2.580 3.700 3.480 ;
        RECT  4.930 2.680 5.210 3.480 ;
        RECT  6.020 2.680 6.300 3.480 ;
        RECT  7.340 2.680 7.620 3.480 ;
        RECT  8.420 2.620 8.700 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  1.020 2.680 1.300 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.580 2.530 3.380 2.690 ;
        RECT  3.220 2.260 3.380 2.690 ;
        RECT  2.580 2.360 2.740 2.690 ;
        RECT  3.860 2.360 7.620 2.520 ;
        RECT  7.460 1.720 7.620 2.520 ;
        RECT  0.160 2.360 2.740 2.520 ;
        RECT  3.220 2.260 4.020 2.420 ;
        RECT  0.160 1.020 0.320 2.520 ;
        RECT  7.460 1.720 8.260 1.880 ;
        RECT  8.100 1.340 8.260 1.880 ;
        RECT  0.160 1.020 0.940 1.180 ;
        RECT  6.960 1.400 7.120 2.160 ;
        RECT  6.640 1.400 7.720 1.560 ;
        RECT  6.640 0.880 6.800 1.560 ;
        RECT  5.480 0.820 5.640 2.160 ;
        RECT  4.860 0.820 6.400 0.980 ;
        RECT  6.240 0.560 6.400 0.980 ;
        RECT  6.240 0.560 6.520 0.720 ;
        RECT  4.180 0.820 4.340 2.160 ;
        RECT  4.180 0.820 4.660 0.980 ;
        RECT  4.500 0.440 4.660 0.980 ;
        RECT  4.500 0.440 4.840 0.600 ;
        RECT  2.900 1.820 3.060 2.320 ;
        RECT  2.920 0.820 3.080 1.980 ;
        RECT  2.580 0.820 3.080 0.980 ;
        RECT  2.640 0.440 2.800 0.980 ;
        RECT  2.400 0.440 2.800 0.600 ;
        RECT  0.860 2.040 1.900 2.200 ;
        RECT  0.860 1.460 1.020 2.200 ;
        RECT  0.860 1.460 1.260 1.620 ;
        RECT  1.100 0.820 1.260 1.620 ;
        RECT  1.100 0.820 2.380 0.980 ;
    END
END ND8DHD

MACRO NR2BHD
    CLASS CORE ;
    FOREIGN NR2BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.680 1.500 2.440 ;
        RECT  1.280 2.160 1.500 2.440 ;
        RECT  0.660 0.680 1.500 0.880 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.040 1.100 1.580 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.420 0.300 1.960 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.400 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
END NR2BHD

MACRO NR2CHD
    CLASS CORE ;
    FOREIGN NR2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.280 2.080 1.500 2.360 ;
        RECT  1.300 0.920 1.500 2.460 ;
        RECT  0.620 0.920 1.500 1.080 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.100 2.000 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 1.130 0.300 1.670 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.760 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
END NR2CHD

MACRO NR2EHD
    CLASS CORE ;
    FOREIGN NR2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.580 2.700 2.280 ;
        RECT  0.100 2.120 2.700 2.280 ;
        RECT  0.100 0.580 2.700 0.780 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.320 1.620 ;
        RECT  0.100 0.940 2.320 1.140 ;
        RECT  2.160 0.940 2.320 1.460 ;
        RECT  0.100 0.940 0.300 1.670 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.420 1.900 1.960 ;
        RECT  1.680 1.460 1.900 1.740 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.060 2.440 1.700 3.480 ;
        END
    END VCC
END NR2EHD

MACRO NR2GHD
    CLASS CORE ;
    FOREIGN NR2GHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.600 3.500 2.440 ;
        RECT  0.100 2.280 3.500 2.440 ;
        RECT  0.540 0.600 3.500 0.760 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.100 0.320 1.620 ;
        RECT  0.100 1.100 2.220 1.300 ;
        RECT  2.060 1.100 2.220 1.440 ;
        RECT  0.100 1.100 0.300 1.960 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.700 3.100 1.900 ;
        RECT  2.900 1.060 3.100 2.070 ;
        RECT  0.900 1.460 1.100 1.900 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.220 -0.280 2.500 0.400 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  1.100 -0.280 1.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.220 2.600 3.500 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  1.060 2.620 1.340 3.480 ;
        END
    END VCC
END NR2GHD

MACRO NR2IHD
    CLASS CORE ;
    FOREIGN NR2IHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.420 2.280 5.100 2.440 ;
        RECT  4.900 0.440 5.100 2.760 ;
        RECT  0.860 0.560 5.100 0.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.380 1.460 3.540 1.900 ;
        RECT  4.500 1.140 4.700 1.900 ;
        RECT  1.700 1.700 4.700 1.900 ;
        RECT  1.700 1.260 1.900 1.970 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.700 0.900 2.860 1.420 ;
        RECT  0.500 0.900 4.020 1.100 ;
        RECT  3.860 0.900 4.020 1.420 ;
        RECT  0.500 0.700 0.700 1.960 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.660 -0.280 3.940 0.400 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  1.420 -0.280 1.700 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 2.620 2.580 3.480 ;
        RECT  3.980 2.600 4.260 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.620 2.440 0.900 3.480 ;
        END
    END VCC
END NR2IHD

MACRO NR3BHD
    CLASS CORE ;
    FOREIGN NR3BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.640 2.300 2.440 ;
        RECT  1.700 2.240 2.300 2.440 ;
        RECT  0.260 0.640 2.300 0.840 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.040 1.140 1.320 ;
        RECT  0.900 1.040 1.100 1.560 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.460 0.700 1.980 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 1.900 1.980 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.940 -0.280 2.220 0.400 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.820 -0.280 1.100 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.540 2.440 0.820 3.480 ;
        END
    END VCC
END NR3BHD

MACRO NR3EHD
    CLASS CORE ;
    FOREIGN NR3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.660 3.500 2.480 ;
        RECT  3.280 2.200 3.500 2.480 ;
        RECT  3.280 0.660 3.500 0.940 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.140 1.100 1.660 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.460 0.300 1.980 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.460 1.500 1.980 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.540 -0.280 1.820 0.400 ;
        RECT  2.700 -0.280 2.980 0.580 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.700 2.440 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.260 2.440 0.540 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.140 1.940 3.080 2.100 ;
        RECT  2.920 0.800 3.080 2.100 ;
        RECT  2.140 0.800 3.080 0.960 ;
        RECT  1.420 2.260 1.880 2.420 ;
        RECT  1.720 0.800 1.880 2.420 ;
        RECT  1.720 1.460 2.600 1.620 ;
        RECT  0.100 0.800 1.880 0.960 ;
        RECT  0.100 0.740 0.380 0.960 ;
    END
END NR3EHD

MACRO NR3HHD
    CLASS CORE ;
    FOREIGN NR3HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.700 3.500 2.500 ;
        RECT  3.090 2.340 3.500 2.500 ;
        RECT  3.090 0.700 3.500 0.860 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.140 1.100 1.660 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.460 0.320 1.740 ;
        RECT  0.100 1.460 0.300 1.980 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.460 1.500 1.980 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.540 -0.280 1.820 0.400 ;
        RECT  2.570 -0.280 2.850 0.860 ;
        RECT  3.680 -0.280 3.900 0.920 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.570 2.340 2.850 3.480 ;
        RECT  3.680 2.280 3.900 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.260 2.440 0.540 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.050 2.020 3.080 2.180 ;
        RECT  2.920 1.020 3.080 2.180 ;
        RECT  2.050 1.020 3.080 1.180 ;
        RECT  1.420 2.260 1.880 2.420 ;
        RECT  1.720 0.800 1.880 2.420 ;
        RECT  1.720 1.460 2.510 1.620 ;
        RECT  0.100 0.800 1.880 0.960 ;
        RECT  0.100 0.740 0.380 0.960 ;
    END
END NR3HHD

MACRO NR4CHD
    CLASS CORE ;
    FOREIGN NR4CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.780 4.300 2.390 ;
        RECT  4.080 2.110 4.300 2.390 ;
        RECT  4.080 0.780 4.300 1.060 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.580 1.500 2.100 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.760 ;
        RECT  2.080 1.240 2.300 1.520 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.840 1.240 1.100 1.520 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.680 0.320 1.960 ;
        RECT  0.100 1.640 0.300 2.160 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 -0.280 1.320 0.400 ;
        RECT  1.980 -0.280 2.260 0.400 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.260 2.440 2.540 3.480 ;
        RECT  3.340 2.800 3.620 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.380 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.780 2.440 3.880 2.600 ;
        RECT  3.720 0.560 3.880 2.600 ;
        RECT  2.460 0.560 3.880 0.720 ;
        RECT  0.940 2.260 1.220 2.480 ;
        RECT  0.520 2.260 1.220 2.420 ;
        RECT  0.520 0.880 0.680 2.420 ;
        RECT  3.120 0.920 3.400 1.110 ;
        RECT  2.120 0.920 3.400 1.080 ;
        RECT  0.660 0.560 0.820 1.040 ;
        RECT  2.120 0.560 2.280 1.080 ;
        RECT  0.660 0.560 2.280 0.720 ;
        RECT  1.420 2.260 1.700 2.480 ;
        RECT  1.420 2.260 1.880 2.420 ;
        RECT  1.720 0.880 1.880 2.420 ;
        RECT  2.500 2.020 2.780 2.280 ;
        RECT  1.720 2.120 2.780 2.280 ;
        RECT  1.540 0.880 1.880 1.100 ;
    END
END NR4CHD

MACRO NR4EHD
    CLASS CORE ;
    FOREIGN NR4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.640 4.300 2.560 ;
        RECT  4.080 2.280 4.300 2.560 ;
        RECT  4.080 0.640 4.300 0.920 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.580 1.500 2.100 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.760 ;
        RECT  2.080 1.240 2.300 1.520 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.840 1.240 1.100 1.520 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.680 0.320 1.960 ;
        RECT  0.100 1.640 0.300 2.160 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 -0.280 1.320 0.400 ;
        RECT  1.980 -0.280 2.260 0.400 ;
        RECT  3.390 -0.280 3.670 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.260 2.440 2.540 3.480 ;
        RECT  3.400 2.800 3.680 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.380 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.780 2.440 3.880 2.600 ;
        RECT  3.720 0.560 3.880 2.600 ;
        RECT  2.460 0.560 3.880 0.720 ;
        RECT  0.940 2.260 1.220 2.480 ;
        RECT  0.520 2.260 1.220 2.420 ;
        RECT  0.520 0.880 0.680 2.420 ;
        RECT  3.120 0.920 3.400 1.110 ;
        RECT  2.120 0.920 3.400 1.080 ;
        RECT  0.660 0.560 0.820 1.040 ;
        RECT  2.120 0.560 2.280 1.080 ;
        RECT  0.660 0.560 2.280 0.720 ;
        RECT  1.420 2.260 1.700 2.480 ;
        RECT  1.420 2.260 1.880 2.420 ;
        RECT  1.720 0.880 1.880 2.420 ;
        RECT  2.500 2.020 2.780 2.280 ;
        RECT  1.720 2.120 2.780 2.280 ;
        RECT  1.540 0.880 1.880 1.100 ;
    END
END NR4EHD

MACRO NR4HHD
    CLASS CORE ;
    FOREIGN NR4HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.640 4.300 2.560 ;
        RECT  3.960 2.280 4.300 2.560 ;
        RECT  3.960 0.640 4.300 0.920 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.580 1.500 2.100 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.760 ;
        RECT  2.040 1.240 2.300 1.520 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.840 1.240 1.100 1.520 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.680 0.320 1.960 ;
        RECT  0.100 1.640 0.300 2.160 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.040 -0.280 1.320 0.400 ;
        RECT  1.980 -0.280 2.260 0.400 ;
        RECT  3.340 -0.280 3.620 0.400 ;
        RECT  4.480 -0.280 4.700 0.640 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.260 2.440 2.540 3.480 ;
        RECT  3.340 2.800 3.620 3.480 ;
        RECT  4.480 2.560 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.380 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.780 2.440 3.660 2.600 ;
        RECT  3.500 0.560 3.660 2.600 ;
        RECT  2.460 0.560 3.660 0.720 ;
        RECT  0.940 2.260 1.220 2.480 ;
        RECT  0.520 2.260 1.220 2.420 ;
        RECT  0.520 0.880 0.680 2.420 ;
        RECT  3.000 0.880 3.160 1.710 ;
        RECT  2.120 0.880 3.160 1.040 ;
        RECT  0.660 0.560 0.820 1.040 ;
        RECT  2.120 0.560 2.280 1.040 ;
        RECT  0.660 0.560 2.280 0.720 ;
        RECT  1.420 2.260 1.700 2.480 ;
        RECT  1.420 2.260 1.880 2.420 ;
        RECT  1.720 0.880 1.880 2.420 ;
        RECT  2.520 1.630 2.680 2.280 ;
        RECT  1.720 2.120 2.680 2.280 ;
        RECT  1.540 0.880 1.880 1.100 ;
    END
END NR4HHD

MACRO NR5EHD
    CLASS CORE ;
    FOREIGN NR5EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.880 0.600 5.080 2.680 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.760 ;
        END
    END I1
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.200 2.700 1.720 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.980 1.240 2.300 1.750 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.800 -0.280 1.960 0.840 ;
        RECT  2.820 -0.280 4.540 0.400 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.320 2.560 3.480 3.480 ;
        RECT  4.360 2.560 4.520 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  1.560 2.800 1.840 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.780 2.600 4.060 2.760 ;
        RECT  3.900 2.220 4.060 2.760 ;
        RECT  3.900 2.220 4.700 2.380 ;
        RECT  4.540 1.390 4.700 2.380 ;
        RECT  3.520 1.390 4.700 1.550 ;
        RECT  3.520 0.880 3.680 1.550 ;
        RECT  2.580 1.880 2.900 2.060 ;
        RECT  2.580 1.880 4.180 2.040 ;
        RECT  4.020 1.760 4.180 2.040 ;
        RECT  3.180 0.620 3.340 2.040 ;
        RECT  2.260 0.620 3.340 0.780 ;
        RECT  0.140 2.420 3.160 2.580 ;
        RECT  3.000 2.240 3.160 2.580 ;
        RECT  0.520 0.620 0.680 2.580 ;
        RECT  3.000 2.240 3.700 2.400 ;
        RECT  3.380 2.200 3.700 2.400 ;
        RECT  0.100 0.620 1.500 0.780 ;
    END
END NR5EHD

MACRO NR6EHD
    CLASS CORE ;
    FOREIGN NR6EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.280 0.600 5.480 2.680 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.230 1.500 1.760 ;
        END
    END I1
    PIN I6
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.160 3.140 1.440 ;
        RECT  2.900 1.160 3.100 1.680 ;
        END
    END I6
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.140 2.700 1.720 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.980 1.240 2.300 1.760 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.800 -0.280 1.960 0.840 ;
        RECT  2.820 -0.280 3.100 0.400 ;
        RECT  4.660 -0.280 4.940 0.400 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.660 2.580 3.940 3.480 ;
        RECT  4.760 2.560 4.920 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  1.610 2.560 1.890 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.180 2.540 4.480 2.760 ;
        RECT  4.320 2.220 4.480 2.760 ;
        RECT  4.320 2.220 5.100 2.380 ;
        RECT  4.940 1.390 5.100 2.380 ;
        RECT  3.920 1.390 5.100 1.550 ;
        RECT  3.920 0.880 4.080 1.550 ;
        RECT  3.060 1.840 3.380 2.060 ;
        RECT  4.420 1.760 4.580 2.040 ;
        RECT  3.060 1.840 4.580 2.000 ;
        RECT  3.540 0.500 3.700 2.000 ;
        RECT  2.260 0.620 3.700 0.780 ;
        RECT  3.420 0.500 3.700 0.780 ;
        RECT  0.140 2.220 4.160 2.380 ;
        RECT  3.840 2.160 4.160 2.380 ;
        RECT  0.520 0.620 0.680 2.380 ;
        RECT  0.100 0.620 1.500 0.780 ;
    END
END NR6EHD

MACRO NR8EHD
    CLASS CORE ;
    FOREIGN NR8EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.800 9.100 2.400 ;
        RECT  7.860 2.200 9.100 2.400 ;
        RECT  8.260 0.800 9.100 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.520 1.520 ;
        RECT  1.300 1.240 1.500 1.760 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.240 0.320 1.520 ;
        RECT  0.100 1.240 0.300 1.760 ;
        END
    END I1
    PIN I8
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 1.240 4.700 1.760 ;
        END
    END I8
    PIN I7
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 1.200 5.900 1.740 ;
        END
    END I7
    PIN I6
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.200 5.260 1.480 ;
        RECT  4.900 1.200 5.100 1.760 ;
        END
    END I6
    PIN I5
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.240 3.980 1.520 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END I5
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.760 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.210 2.040 1.490 ;
        RECT  1.700 1.210 1.900 1.730 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.200 -0.280 1.360 0.840 ;
        RECT  2.220 -0.280 2.500 0.400 ;
        RECT  3.740 -0.280 6.320 0.400 ;
        RECT  7.410 -0.280 7.690 0.400 ;
        RECT  8.820 -0.280 9.040 0.640 ;
        RECT  0.000 -0.280 9.200 0.280 ;
        RECT  0.160 -0.280 0.320 0.840 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.440 2.560 2.600 3.480 ;
        RECT  3.480 2.560 3.640 3.480 ;
        RECT  4.660 2.800 4.940 3.480 ;
        RECT  6.040 2.560 6.200 3.480 ;
        RECT  7.080 2.560 7.300 3.480 ;
        RECT  8.820 2.560 9.040 3.480 ;
        RECT  0.000 2.920 9.200 3.480 ;
        RECT  1.020 2.800 1.300 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.500 2.600 6.920 2.760 ;
        RECT  6.760 2.220 6.920 2.760 ;
        RECT  6.760 2.220 7.460 2.380 ;
        RECT  7.300 0.920 7.460 2.380 ;
        RECT  7.300 1.830 8.740 1.990 ;
        RECT  8.580 1.390 8.740 1.990 ;
        RECT  7.260 1.390 7.460 1.670 ;
        RECT  2.900 2.600 3.180 2.760 ;
        RECT  3.020 2.220 3.180 2.760 ;
        RECT  3.020 2.220 3.540 2.380 ;
        RECT  3.380 0.560 3.540 2.380 ;
        RECT  7.870 0.560 8.030 1.670 ;
        RECT  2.640 0.560 2.800 1.100 ;
        RECT  2.640 0.560 8.030 0.720 ;
        RECT  4.180 2.240 6.600 2.400 ;
        RECT  6.440 1.900 6.600 2.400 ;
        RECT  4.180 0.880 4.340 2.400 ;
        RECT  3.740 1.990 4.340 2.150 ;
        RECT  6.440 1.900 6.960 2.060 ;
        RECT  4.180 0.880 4.620 1.040 ;
        RECT  5.900 1.920 6.260 2.080 ;
        RECT  6.100 0.880 6.260 2.080 ;
        RECT  6.100 1.400 6.650 1.560 ;
        RECT  5.440 0.880 6.260 1.040 ;
        RECT  1.980 1.920 2.400 2.080 ;
        RECT  2.240 0.620 2.400 2.080 ;
        RECT  2.240 1.600 3.220 1.760 ;
        RECT  1.660 0.620 2.400 0.780 ;
        RECT  0.100 2.240 2.840 2.400 ;
        RECT  2.560 2.120 2.840 2.400 ;
        RECT  0.520 0.620 0.680 2.400 ;
        RECT  0.520 0.620 0.900 0.780 ;
    END
END NR8EHD

MACRO OA112CHD
    CLASS CORE ;
    FOREIGN OA112CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.600 0.960 2.760 1.240 ;
        RECT  2.600 1.040 3.100 1.240 ;
        RECT  2.900 1.040 3.100 2.440 ;
        RECT  2.570 2.240 3.100 2.440 ;
        RECT  2.570 2.240 2.730 2.520 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.510 1.520 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.210 -0.280 3.490 0.820 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.030 2.620 3.310 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.480 2.470 1.760 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
    END
END OA112CHD

MACRO OA112EHD
    CLASS CORE ;
    FOREIGN OA112EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.700 1.010 3.100 1.210 ;
        RECT  2.900 1.010 3.100 2.440 ;
        RECT  2.570 2.240 3.100 2.440 ;
        RECT  2.570 2.240 2.730 2.520 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.260 1.510 1.540 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.220 -0.280 3.500 0.820 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.030 2.620 3.310 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.460 2.470 1.740 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
    END
END OA112EHD

MACRO OA112HHD
    CLASS CORE ;
    FOREIGN OA112HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.920 3.500 2.420 ;
        RECT  2.570 2.260 3.900 2.420 ;
        RECT  2.700 0.920 4.090 1.080 ;
        RECT  2.570 2.240 2.730 2.520 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.260 1.510 1.540 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.220 -0.280 3.500 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.030 2.620 3.310 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.460 2.470 1.740 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
    END
END OA112HHD

MACRO OA112KHD
    CLASS CORE ;
    FOREIGN OA112KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.920 3.900 2.420 ;
        RECT  2.570 2.260 4.970 2.420 ;
        RECT  4.810 0.860 5.090 1.080 ;
        RECT  2.700 0.920 5.090 1.080 ;
        RECT  2.570 2.240 2.730 2.520 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.260 1.510 1.540 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.220 -0.280 3.500 0.580 ;
        RECT  4.260 -0.280 4.540 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.030 2.620 3.310 3.480 ;
        RECT  4.100 2.620 4.380 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.460 2.470 1.740 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
    END
END OA112KHD

MACRO OA12CHD
    CLASS CORE ;
    FOREIGN OA12CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.000 2.700 2.460 ;
        RECT  2.230 2.260 2.700 2.460 ;
        RECT  2.260 1.000 2.700 1.200 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.200 1.100 1.800 ;
        RECT  0.860 1.200 1.100 1.480 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.520 1.510 1.800 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.820 -0.280 3.100 0.820 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  1.780 -0.280 2.060 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.560 2.320 1.720 3.480 ;
        RECT  1.560 2.320 1.780 2.600 ;
        RECT  2.750 2.620 3.030 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.370 2.580 ;
        RECT  1.210 2.000 1.370 2.580 ;
        RECT  1.210 2.000 2.020 2.160 ;
        RECT  1.720 1.860 2.020 2.160 ;
        RECT  1.720 0.760 1.880 2.160 ;
        RECT  0.640 0.760 1.880 0.920 ;
        RECT  0.100 0.440 0.380 0.660 ;
        RECT  0.100 0.440 1.580 0.600 ;
    END
END OA12CHD

MACRO OA12EHD
    CLASS CORE ;
    FOREIGN OA12EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.900 2.700 2.460 ;
        RECT  2.230 2.260 2.700 2.460 ;
        RECT  2.260 0.900 2.700 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.860 1.520 1.100 1.800 ;
        RECT  0.900 1.200 1.100 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.720 1.600 1.880 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.820 -0.280 3.100 0.580 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  1.780 -0.280 2.060 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  2.750 2.620 3.030 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.060 1.340 2.580 ;
        RECT  1.180 2.060 2.050 2.220 ;
        RECT  1.890 0.760 2.050 2.220 ;
        RECT  0.680 0.760 2.050 0.920 ;
        RECT  0.160 0.440 0.320 1.000 ;
        RECT  0.160 0.440 1.580 0.600 ;
    END
END OA12EHD

MACRO OA12HHD
    CLASS CORE ;
    FOREIGN OA12HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.540 0.860 2.820 1.080 ;
        RECT  2.540 0.920 3.900 1.080 ;
        RECT  3.300 0.920 3.500 2.460 ;
        RECT  2.510 2.300 3.870 2.460 ;
        RECT  3.300 0.920 3.900 1.140 ;
        RECT  2.510 2.300 2.790 2.520 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.100 2.040 ;
        RECT  0.860 1.460 1.100 1.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.660 1.590 1.940 ;
        RECT  1.300 1.400 1.500 2.040 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 -0.280 3.380 0.580 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  1.780 -0.280 2.060 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.520 1.780 3.480 ;
        RECT  3.030 2.620 3.310 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.200 1.340 2.580 ;
        RECT  1.180 2.200 2.350 2.360 ;
        RECT  2.190 0.940 2.350 2.360 ;
        RECT  0.640 0.940 2.350 1.100 ;
        RECT  0.100 0.620 1.540 0.780 ;
    END
END OA12HHD

MACRO OA12KHD
    CLASS CORE ;
    FOREIGN OA12KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.300 5.070 2.460 ;
        RECT  4.820 0.860 5.100 1.080 ;
        RECT  2.740 0.920 5.100 1.080 ;
        RECT  3.700 0.920 3.900 2.460 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.100 2.040 ;
        RECT  0.860 1.460 1.100 1.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.660 1.590 1.940 ;
        RECT  1.300 1.400 1.500 2.040 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.260 -0.280 3.540 0.580 ;
        RECT  4.300 -0.280 4.580 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  1.780 -0.280 2.060 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.620 1.780 3.480 ;
        RECT  3.150 2.620 3.430 3.480 ;
        RECT  4.230 2.620 4.510 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.300 2.350 2.460 ;
        RECT  2.190 0.940 2.350 2.460 ;
        RECT  0.640 0.940 2.350 1.100 ;
        RECT  0.100 0.620 1.540 0.780 ;
    END
END OA12KHD

MACRO OA13CHD
    CLASS CORE ;
    FOREIGN OA13CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.660 3.100 2.640 ;
        RECT  2.830 2.360 3.100 2.640 ;
        RECT  2.880 0.660 3.100 0.940 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.080 1.240 2.300 1.520 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        RECT  1.540 1.240 1.900 1.520 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.180 1.580 ;
        RECT  0.900 1.240 1.100 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.490 1.300 0.700 1.580 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 -0.280 2.580 0.810 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  1.140 -0.280 1.420 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.120 2.430 0.400 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 2.600 2.020 2.760 ;
        RECT  1.860 2.300 2.020 2.760 ;
        RECT  0.560 2.110 0.720 2.760 ;
        RECT  1.860 2.300 2.670 2.460 ;
        RECT  2.510 1.620 2.670 2.460 ;
        RECT  0.160 2.110 0.720 2.270 ;
        RECT  0.160 0.660 0.320 2.270 ;
        RECT  0.680 0.920 1.880 1.080 ;
        RECT  1.720 0.660 1.880 1.080 ;
        RECT  0.680 0.660 0.840 1.080 ;
    END
END OA13CHD

MACRO OA13EHD
    CLASS CORE ;
    FOREIGN OA13EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.660 3.100 2.640 ;
        RECT  2.830 2.360 3.100 2.640 ;
        RECT  2.880 0.660 3.100 0.940 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.060 1.240 2.300 1.520 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        RECT  1.540 1.240 1.900 1.520 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.300 1.180 1.580 ;
        RECT  0.900 1.240 1.100 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.490 1.340 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 -0.280 2.580 0.810 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  1.220 -0.280 1.500 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.120 2.430 0.400 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 2.600 2.020 2.760 ;
        RECT  1.860 2.300 2.020 2.760 ;
        RECT  0.560 2.110 0.720 2.760 ;
        RECT  1.860 2.300 2.670 2.460 ;
        RECT  2.510 1.460 2.670 2.460 ;
        RECT  0.160 2.110 0.720 2.270 ;
        RECT  0.160 0.660 0.320 2.270 ;
        RECT  2.510 1.460 2.700 1.740 ;
        RECT  0.700 0.920 1.960 1.080 ;
        RECT  1.800 0.660 1.960 1.080 ;
    END
END OA13EHD

MACRO OA13HHD
    CLASS CORE ;
    FOREIGN OA13HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.840 3.100 2.760 ;
        RECT  2.620 2.600 3.100 2.760 ;
        RECT  2.760 0.840 3.100 1.120 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.060 1.460 2.300 1.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        RECT  1.540 1.460 1.900 1.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.180 1.740 ;
        RECT  0.900 1.240 1.100 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.490 1.340 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 -0.280 2.460 0.580 ;
        RECT  3.220 -0.280 3.500 0.660 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  1.140 -0.280 1.420 0.660 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.140 2.620 2.420 3.480 ;
        RECT  3.280 2.520 3.440 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.120 2.410 0.400 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 2.600 1.980 2.760 ;
        RECT  1.820 2.280 1.980 2.760 ;
        RECT  0.560 2.090 0.720 2.760 ;
        RECT  1.820 2.280 2.670 2.440 ;
        RECT  2.510 1.460 2.670 2.440 ;
        RECT  0.160 2.090 0.720 2.250 ;
        RECT  0.160 0.620 0.320 2.250 ;
        RECT  2.510 1.460 2.700 1.740 ;
        RECT  0.620 0.820 1.940 0.980 ;
    END
END OA13HHD

MACRO OA13KHD
    CLASS CORE ;
    FOREIGN OA13KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.740 3.500 2.280 ;
        RECT  2.700 0.740 4.060 0.900 ;
        RECT  2.830 2.120 4.170 2.280 ;
        RECT  2.830 2.060 2.990 2.340 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.060 1.460 2.300 1.740 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        RECT  1.540 1.460 1.900 1.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.180 1.740 ;
        RECT  0.900 1.240 1.100 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.490 1.340 0.700 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 -0.280 2.460 0.580 ;
        RECT  3.260 -0.280 3.540 0.580 ;
        RECT  4.340 -0.280 4.620 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  1.140 -0.280 1.420 0.660 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 2.620 2.460 3.480 ;
        RECT  3.300 2.620 3.580 3.480 ;
        RECT  4.380 2.620 4.660 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.120 2.410 0.400 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.560 2.600 2.020 2.760 ;
        RECT  1.860 2.300 2.020 2.760 ;
        RECT  0.560 2.090 0.720 2.760 ;
        RECT  1.860 2.300 2.670 2.460 ;
        RECT  2.510 1.460 2.670 2.460 ;
        RECT  0.160 2.090 0.720 2.250 ;
        RECT  0.160 0.660 0.320 2.250 ;
        RECT  2.510 1.460 2.700 1.740 ;
        RECT  0.620 0.820 1.940 0.980 ;
    END
END OA13KHD

MACRO OA2222CHD
    CLASS CORE ;
    FOREIGN OA2222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.840 0.540 6.000 1.140 ;
        RECT  5.840 0.980 6.700 1.140 ;
        RECT  6.500 0.980 6.700 2.460 ;
        RECT  5.320 2.300 6.700 2.460 ;
        RECT  5.320 2.300 5.480 2.640 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.240 5.100 1.800 ;
        RECT  4.640 1.340 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.260 -0.280 5.540 0.760 ;
        RECT  6.300 -0.280 6.580 0.760 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.420 2.270 3.480 ;
        RECT  2.660 2.420 2.940 3.480 ;
        RECT  4.540 2.580 4.820 3.480 ;
        RECT  6.300 2.620 6.580 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.100 2.260 5.160 2.420 ;
        RECT  5.000 1.960 5.160 2.420 ;
        RECT  0.940 2.100 3.260 2.260 ;
        RECT  5.000 1.960 6.140 2.120 ;
        RECT  5.980 1.450 6.140 2.120 ;
        RECT  1.720 0.820 1.880 2.260 ;
        RECT  1.660 0.820 1.940 0.980 ;
        RECT  3.500 1.930 4.380 2.090 ;
        RECT  4.220 0.820 4.380 2.090 ;
        RECT  5.450 0.920 5.610 1.570 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  4.220 0.820 4.500 1.080 ;
        RECT  2.720 0.920 3.920 1.080 ;
        RECT  3.760 0.500 3.920 1.080 ;
        RECT  2.720 0.720 2.880 1.080 ;
        RECT  4.740 0.500 5.020 0.760 ;
        RECT  3.760 0.500 5.020 0.660 ;
        RECT  0.100 0.920 1.360 1.080 ;
        RECT  1.200 0.500 1.360 1.080 ;
        RECT  0.160 0.660 0.320 1.080 ;
        RECT  2.180 0.500 2.460 0.760 ;
        RECT  1.200 0.500 2.460 0.660 ;
    END
END OA2222CHD

MACRO OA2222EHD
    CLASS CORE ;
    FOREIGN OA2222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.800 0.500 5.960 1.040 ;
        RECT  5.800 0.880 7.500 1.040 ;
        RECT  7.300 0.880 7.500 2.460 ;
        RECT  5.330 2.300 7.500 2.460 ;
        RECT  5.330 2.300 5.490 2.640 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.240 5.100 1.800 ;
        RECT  4.640 1.340 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.220 -0.280 5.500 0.760 ;
        RECT  6.260 -0.280 6.540 0.720 ;
        RECT  7.300 -0.280 7.580 0.720 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 2.580 2.930 3.480 ;
        RECT  4.550 2.560 4.830 3.480 ;
        RECT  6.110 2.620 6.390 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.500 1.920 4.380 2.080 ;
        RECT  4.220 0.920 4.380 2.080 ;
        RECT  6.980 1.200 7.140 1.660 ;
        RECT  5.450 0.920 5.610 1.620 ;
        RECT  5.450 1.200 7.140 1.360 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  0.940 2.240 5.160 2.400 ;
        RECT  5.000 1.960 5.160 2.400 ;
        RECT  1.720 0.920 1.880 2.400 ;
        RECT  5.000 1.960 6.420 2.120 ;
        RECT  6.200 1.520 6.420 2.120 ;
        RECT  6.200 1.520 6.480 1.680 ;
        RECT  1.660 0.920 1.940 1.080 ;
        RECT  2.620 0.920 3.980 1.080 ;
        RECT  3.820 0.600 3.980 1.080 ;
        RECT  3.820 0.600 5.020 0.760 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OA2222EHD

MACRO OA2222HHD
    CLASS CORE ;
    FOREIGN OA2222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.330 2.110 5.740 2.270 ;
        RECT  5.800 0.500 5.960 1.040 ;
        RECT  5.800 0.880 9.900 1.040 ;
        RECT  5.580 1.970 9.900 2.130 ;
        RECT  9.700 0.880 9.900 2.130 ;
        RECT  5.330 2.110 5.490 2.640 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.640 1.340 5.100 1.620 ;
        RECT  4.900 1.240 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.220 -0.280 5.500 0.760 ;
        RECT  6.260 -0.280 6.540 0.720 ;
        RECT  7.300 -0.280 7.580 0.720 ;
        RECT  8.340 -0.280 8.620 0.720 ;
        RECT  9.390 -0.280 9.670 0.720 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 2.580 2.930 3.480 ;
        RECT  4.550 2.560 4.830 3.480 ;
        RECT  6.310 2.620 6.590 3.480 ;
        RECT  8.410 2.620 8.690 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.500 1.920 4.380 2.080 ;
        RECT  4.220 0.920 4.380 2.080 ;
        RECT  9.130 1.200 9.290 1.620 ;
        RECT  7.110 1.200 7.750 1.480 ;
        RECT  5.390 1.320 5.670 1.480 ;
        RECT  5.450 1.200 9.290 1.360 ;
        RECT  5.450 0.920 5.610 1.480 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  7.890 2.300 9.210 2.460 ;
        RECT  0.940 2.240 5.160 2.400 ;
        RECT  5.000 1.780 5.160 2.400 ;
        RECT  1.720 0.920 1.880 2.400 ;
        RECT  5.000 1.780 5.420 1.940 ;
        RECT  8.280 1.520 8.560 1.800 ;
        RECT  5.260 1.640 8.560 1.800 ;
        RECT  6.200 1.520 6.480 1.800 ;
        RECT  1.660 0.920 1.940 1.080 ;
        RECT  5.790 2.510 6.070 2.670 ;
        RECT  5.910 2.300 6.070 2.670 ;
        RECT  5.910 2.300 7.130 2.460 ;
        RECT  2.620 0.920 3.980 1.080 ;
        RECT  3.820 0.600 3.980 1.080 ;
        RECT  3.820 0.600 5.020 0.760 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OA2222HHD

MACRO OA222CHD
    CLASS CORE ;
    FOREIGN OA222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.240 0.980 4.700 1.140 ;
        RECT  4.500 0.980 4.700 2.280 ;
        RECT  4.040 2.060 4.700 2.280 ;
        RECT  4.240 0.800 4.400 1.140 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.720 ;
        RECT  4.700 -0.280 4.980 0.820 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.620 2.840 3.480 ;
        RECT  4.630 2.440 4.910 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.520 2.300 3.880 2.460 ;
        RECT  3.720 1.470 3.880 2.460 ;
        RECT  3.720 1.470 4.060 1.630 ;
        RECT  3.900 0.880 4.060 1.630 ;
        RECT  3.140 0.880 4.060 1.040 ;
        RECT  1.620 0.560 3.980 0.720 ;
        RECT  0.580 0.880 2.420 1.040 ;
    END
END OA222CHD

MACRO OA222EHD
    CLASS CORE ;
    FOREIGN OA222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.240 0.920 4.700 1.080 ;
        RECT  4.500 0.920 4.700 2.280 ;
        RECT  4.040 2.060 4.700 2.280 ;
        RECT  4.240 0.760 4.400 1.080 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  4.700 -0.280 4.980 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.100 -0.280 0.380 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.620 2.840 3.480 ;
        RECT  4.630 2.620 4.910 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.480 2.260 3.880 2.420 ;
        RECT  3.720 1.470 3.880 2.420 ;
        RECT  3.720 1.470 4.060 1.630 ;
        RECT  3.900 0.760 4.060 1.630 ;
        RECT  3.140 0.760 4.060 0.920 ;
        RECT  1.580 0.440 4.020 0.600 ;
        RECT  0.620 0.760 2.420 0.920 ;
    END
END OA222EHD

MACRO OA222HHD
    CLASS CORE ;
    FOREIGN OA222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.240 0.760 4.400 1.080 ;
        RECT  4.900 0.920 5.100 2.280 ;
        RECT  5.220 0.860 5.500 1.080 ;
        RECT  4.240 0.920 5.500 1.080 ;
        RECT  4.040 2.120 5.500 2.280 ;
        RECT  4.040 2.060 4.320 2.280 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  4.700 -0.280 4.980 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.620 2.840 3.480 ;
        RECT  4.630 2.620 4.910 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.480 2.260 3.880 2.420 ;
        RECT  3.720 1.470 3.880 2.420 ;
        RECT  3.720 1.470 4.060 1.630 ;
        RECT  3.900 0.760 4.060 1.630 ;
        RECT  3.140 0.760 4.060 0.920 ;
        RECT  1.580 0.440 4.020 0.600 ;
        RECT  0.620 0.760 2.420 0.920 ;
    END
END OA222HHD

MACRO OA222KHD
    CLASS CORE ;
    FOREIGN OA222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.240 0.760 4.400 1.080 ;
        RECT  4.900 0.920 5.100 2.280 ;
        RECT  4.240 0.920 6.640 1.080 ;
        RECT  4.040 2.120 6.640 2.280 ;
        RECT  4.040 2.060 4.320 2.280 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.580 ;
        RECT  4.700 -0.280 4.980 0.580 ;
        RECT  5.740 -0.280 6.020 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.860 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.620 2.840 3.480 ;
        RECT  4.630 2.620 4.910 3.480 ;
        RECT  5.770 2.620 6.050 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.480 2.260 3.880 2.420 ;
        RECT  3.720 1.470 3.880 2.420 ;
        RECT  3.720 1.470 4.060 1.630 ;
        RECT  3.900 0.760 4.060 1.630 ;
        RECT  3.140 0.760 4.060 0.920 ;
        RECT  1.580 0.440 4.020 0.600 ;
        RECT  0.620 0.760 2.420 0.920 ;
    END
END OA222KHD

MACRO OA22CHD
    CLASS CORE ;
    FOREIGN OA22CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.720 3.100 2.120 ;
        RECT  2.720 1.840 3.100 2.120 ;
        RECT  2.760 0.720 3.100 1.000 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.020 1.620 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.280 -0.280 3.440 1.040 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.440 2.270 3.480 ;
        RECT  3.280 2.120 3.440 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.120 2.550 2.280 ;
        RECT  2.390 0.820 2.550 2.280 ;
        RECT  1.660 0.820 2.550 0.980 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.500 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
        RECT  1.260 0.500 2.540 0.660 ;
    END
END OA22CHD

MACRO OA22EHD
    CLASS CORE ;
    FOREIGN OA22EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.720 3.100 2.340 ;
        RECT  2.720 2.060 3.100 2.340 ;
        RECT  2.720 0.720 3.100 1.000 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.020 1.620 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.280 -0.280 3.440 1.040 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.440 2.270 3.480 ;
        RECT  3.280 2.120 3.440 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.440 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.120 2.550 2.280 ;
        RECT  2.390 0.920 2.550 2.280 ;
        RECT  1.620 0.920 2.550 1.080 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OA22EHD

MACRO OA22HHD
    CLASS CORE ;
    FOREIGN OA22HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.030 2.060 3.250 2.340 ;
        RECT  2.970 0.920 4.300 1.080 ;
        RECT  3.700 0.920 3.900 2.280 ;
        RECT  3.700 0.920 4.300 1.140 ;
        RECT  3.700 2.060 4.300 2.280 ;
        RECT  3.030 2.120 4.300 2.280 ;
        RECT  2.970 0.860 3.250 1.080 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.020 1.620 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.490 -0.280 3.770 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.970 2.620 2.250 3.480 ;
        RECT  3.490 2.620 3.770 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.300 2.810 2.460 ;
        RECT  2.650 0.920 2.810 2.460 ;
        RECT  1.660 0.920 2.810 1.080 ;
        RECT  0.100 0.740 1.420 0.900 ;
        RECT  1.260 0.440 1.420 0.900 ;
        RECT  2.180 0.440 2.460 0.760 ;
        RECT  1.260 0.440 2.460 0.600 ;
    END
END OA22HHD

MACRO OA22KHD
    CLASS CORE ;
    FOREIGN OA22KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.030 2.060 3.250 2.340 ;
        RECT  4.100 0.920 4.300 2.280 ;
        RECT  2.970 0.920 5.390 1.080 ;
        RECT  3.030 2.120 5.390 2.280 ;
        RECT  2.970 0.860 3.250 1.080 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.340 2.020 1.620 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.490 -0.280 3.770 0.580 ;
        RECT  4.540 -0.280 4.820 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.970 2.620 2.250 3.480 ;
        RECT  3.490 2.620 3.770 3.480 ;
        RECT  4.540 2.620 4.820 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.940 2.300 2.810 2.460 ;
        RECT  2.650 0.920 2.810 2.460 ;
        RECT  1.660 0.920 2.810 1.080 ;
        RECT  0.100 0.740 1.420 0.900 ;
        RECT  1.260 0.440 1.420 0.900 ;
        RECT  2.180 0.440 2.460 0.760 ;
        RECT  1.260 0.440 2.460 0.600 ;
    END
END OA22KHD

MACRO OAI112BHD
    CLASS CORE ;
    FOREIGN OAI112BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  2.480 0.740 2.700 1.020 ;
        RECT  1.180 2.000 2.700 2.160 ;
        RECT  2.500 0.740 2.700 2.600 ;
        RECT  2.480 2.320 2.700 2.600 ;
        RECT  1.180 2.000 1.340 2.580 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.510 1.520 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 0.920 1.460 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
    END
END OAI112BHD

MACRO OAI112EHD
    CLASS CORE ;
    FOREIGN OAI112EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.900 3.900 2.300 ;
        RECT  3.550 2.100 3.900 2.300 ;
        RECT  3.580 0.900 3.900 1.100 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.510 1.520 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.060 -0.280 3.340 1.110 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.030 2.620 3.310 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.570 2.360 2.790 2.640 ;
        RECT  2.630 0.930 2.790 2.640 ;
        RECT  3.240 1.420 3.520 1.640 ;
        RECT  2.630 1.420 3.520 1.580 ;
        RECT  2.600 0.930 2.790 1.210 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.480 2.470 1.760 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
    END
END OAI112EHD

MACRO OAI112HHD
    CLASS CORE ;
    FOREIGN OAI112HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.650 2.100 4.300 2.300 ;
        RECT  3.650 0.900 4.300 1.100 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.510 1.520 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.090 -0.280 3.370 0.860 ;
        RECT  4.170 -0.280 4.450 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.080 2.620 3.360 3.480 ;
        RECT  4.190 2.620 4.470 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.620 2.140 2.810 2.420 ;
        RECT  2.650 0.840 2.810 2.420 ;
        RECT  2.650 1.420 3.750 1.580 ;
        RECT  2.630 0.880 2.810 1.160 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.480 2.470 1.760 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.460 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
    END
END OAI112HHD

MACRO OAI112KHD
    CLASS CORE ;
    FOREIGN OAI112KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.620 0.900 4.960 1.100 ;
        RECT  3.620 2.100 4.960 2.300 ;
        RECT  4.100 0.900 4.300 2.300 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.510 1.520 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.520 1.990 1.800 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.820 1.300 1.100 1.580 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.100 -0.280 3.380 0.580 ;
        RECT  4.140 -0.280 4.420 0.580 ;
        RECT  5.200 -0.280 5.480 0.580 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.380 1.780 3.480 ;
        RECT  3.100 2.620 3.380 3.480 ;
        RECT  4.160 2.620 4.440 3.480 ;
        RECT  5.200 2.620 5.480 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.630 0.880 2.790 2.380 ;
        RECT  2.630 2.060 2.800 2.340 ;
        RECT  2.630 1.420 3.940 1.580 ;
        RECT  2.600 0.880 2.790 1.160 ;
        RECT  0.940 2.420 1.340 2.580 ;
        RECT  1.180 2.000 1.340 2.580 ;
        RECT  2.020 2.380 2.410 2.540 ;
        RECT  2.250 0.800 2.410 2.540 ;
        RECT  1.180 2.000 2.410 2.160 ;
        RECT  2.250 1.460 2.470 1.740 ;
        RECT  1.940 0.800 2.410 0.960 ;
        RECT  0.100 0.920 1.460 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
    END
END OAI112KHD

MACRO OAI12CHD
    CLASS CORE ;
    FOREIGN OAI12CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.940 2.420 1.370 2.580 ;
        RECT  1.700 0.740 1.900 2.160 ;
        RECT  1.210 2.000 1.900 2.160 ;
        RECT  1.210 2.000 1.370 2.580 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.300 1.100 1.580 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.510 1.580 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.400 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.560 2.320 1.720 3.480 ;
        RECT  1.560 2.320 1.780 2.600 ;
        RECT  0.000 2.920 2.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
    END
END OAI12CHD

MACRO OAI12EHD
    CLASS CORE ;
    FOREIGN OAI12EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 0.880 3.500 2.340 ;
        RECT  3.280 2.060 3.500 2.340 ;
        RECT  3.260 0.880 3.500 1.160 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.300 1.100 1.580 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.510 1.520 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.680 -0.280 2.960 1.060 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.560 2.320 1.720 3.480 ;
        RECT  2.700 2.620 2.980 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.170 2.360 2.360 2.640 ;
        RECT  2.200 0.880 2.360 2.640 ;
        RECT  2.860 1.420 3.140 1.640 ;
        RECT  2.200 1.420 3.140 1.580 ;
        RECT  0.940 2.420 1.370 2.580 ;
        RECT  1.210 2.000 1.370 2.580 ;
        RECT  1.210 2.000 1.900 2.160 ;
        RECT  1.700 0.740 1.900 2.160 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.140 0.820 1.420 1.080 ;
        RECT  0.100 0.820 0.380 1.080 ;
    END
END OAI12EHD

MACRO OAI12HHD
    CLASS CORE ;
    FOREIGN OAI12HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.480 2.100 4.300 2.300 ;
        RECT  3.480 0.900 4.300 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.300 1.100 1.580 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.590 1.580 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.960 -0.280 3.240 0.860 ;
        RECT  4.000 -0.280 4.280 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.460 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 2.320 1.760 3.480 ;
        RECT  1.600 2.320 1.820 2.600 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.450 2.060 2.640 2.340 ;
        RECT  2.480 0.880 2.640 2.340 ;
        RECT  2.480 1.420 3.580 1.580 ;
        RECT  2.460 0.880 2.640 1.160 ;
        RECT  0.940 2.420 1.370 2.580 ;
        RECT  1.210 2.000 1.370 2.580 ;
        RECT  1.210 2.000 2.110 2.160 ;
        RECT  1.950 0.740 2.110 2.160 ;
        RECT  1.800 0.740 2.110 1.020 ;
        RECT  0.100 0.620 1.500 0.780 ;
    END
END OAI12HHD

MACRO OAI12KHD
    CLASS CORE ;
    FOREIGN OAI12KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 0.900 4.580 1.100 ;
        RECT  3.240 2.100 4.580 2.300 ;
        RECT  4.100 0.900 4.300 2.300 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.300 1.100 1.580 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.510 1.580 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.720 -0.280 3.000 0.580 ;
        RECT  3.760 -0.280 4.040 0.580 ;
        RECT  4.820 -0.280 5.100 0.580 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.560 2.320 1.720 3.480 ;
        RECT  1.560 2.320 1.780 2.600 ;
        RECT  2.720 2.620 3.000 3.480 ;
        RECT  3.780 2.620 4.060 3.480 ;
        RECT  4.820 2.620 5.100 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.240 2.060 2.440 2.340 ;
        RECT  2.240 0.880 2.400 2.340 ;
        RECT  2.240 1.420 3.740 1.580 ;
        RECT  0.940 2.420 1.370 2.580 ;
        RECT  1.210 2.000 1.370 2.580 ;
        RECT  1.210 2.000 1.990 2.160 ;
        RECT  1.830 0.740 1.990 2.160 ;
        RECT  1.720 0.740 1.990 1.020 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
    END
END OAI12KHD

MACRO OAI13BHD
    CLASS CORE ;
    FOREIGN OAI13BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.180 0.880 2.700 1.080 ;
        RECT  2.500 0.880 2.700 2.210 ;
        RECT  1.460 2.050 2.700 2.210 ;
        RECT  2.180 0.820 2.460 1.080 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.540 1.580 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.060 1.300 2.300 1.580 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.760 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.090 2.370 2.370 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.620 0.920 1.940 1.080 ;
        RECT  1.660 0.820 1.940 1.080 ;
        RECT  0.620 0.820 0.900 1.080 ;
    END
END OAI13BHD

MACRO OAI13EHD
    CLASS CORE ;
    FOREIGN OAI13EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.700 2.100 4.300 2.300 ;
        RECT  3.730 0.900 4.300 1.100 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.540 1.580 ;
        RECT  1.300 1.240 1.500 1.790 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.300 2.020 1.580 ;
        RECT  1.700 1.240 1.900 1.790 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.760 ;
        RECT  3.210 -0.280 3.490 1.060 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 2.270 2.360 3.480 ;
        RECT  3.180 2.620 3.460 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.470 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.720 2.360 2.910 2.640 ;
        RECT  2.750 0.880 2.910 2.640 ;
        RECT  2.750 1.420 3.690 1.580 ;
        RECT  1.460 1.950 1.740 2.210 ;
        RECT  1.460 1.950 2.540 2.110 ;
        RECT  2.380 0.720 2.540 2.110 ;
        RECT  2.180 0.720 2.540 0.880 ;
        RECT  0.620 0.920 1.940 1.080 ;
        RECT  1.660 0.720 1.940 1.080 ;
        RECT  0.620 0.720 0.900 1.080 ;
    END
END OAI13EHD

MACRO OAI13HHD
    CLASS CORE ;
    FOREIGN OAI13HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.900 4.700 2.300 ;
        RECT  3.880 2.100 4.700 2.300 ;
        RECT  3.880 0.900 4.700 1.100 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.540 1.580 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.040 1.300 2.300 1.580 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.760 ;
        RECT  3.360 -0.280 3.640 0.860 ;
        RECT  4.400 -0.280 4.680 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 2.370 2.360 3.480 ;
        RECT  3.380 2.620 3.660 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.850 2.140 3.040 2.420 ;
        RECT  2.880 0.840 3.040 2.420 ;
        RECT  2.880 1.420 3.980 1.580 ;
        RECT  2.860 0.840 3.080 1.160 ;
        RECT  1.460 2.050 2.680 2.210 ;
        RECT  2.520 0.820 2.680 2.210 ;
        RECT  2.180 0.820 2.680 0.980 ;
        RECT  0.580 0.920 1.980 1.080 ;
    END
END OAI13HHD

MACRO OAI13KHD
    CLASS CORE ;
    FOREIGN OAI13KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 0.900 5.230 1.100 ;
        RECT  3.890 2.100 5.230 2.300 ;
        RECT  4.500 0.900 4.700 2.300 ;
        END
    END O
    PIN B3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B3
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.300 1.540 1.580 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  2.040 1.300 2.300 1.580 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.760 ;
        RECT  3.370 -0.280 3.650 0.580 ;
        RECT  4.410 -0.280 4.690 0.580 ;
        RECT  5.470 -0.280 5.750 0.580 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.080 2.370 2.360 3.480 ;
        RECT  3.370 2.620 3.650 3.480 ;
        RECT  4.430 2.620 4.710 3.480 ;
        RECT  5.470 2.620 5.750 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.890 2.060 3.130 2.380 ;
        RECT  2.890 0.840 3.050 2.380 ;
        RECT  2.890 1.420 4.340 1.580 ;
        RECT  2.870 0.840 3.090 1.160 ;
        RECT  1.460 2.050 2.680 2.210 ;
        RECT  2.520 0.820 2.680 2.210 ;
        RECT  2.180 0.820 2.680 0.980 ;
        RECT  0.580 0.920 1.980 1.080 ;
    END
END OAI13KHD

MACRO OAI2222CHD
    CLASS CORE ;
    FOREIGN OAI2222CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.700 7.100 2.550 ;
        RECT  6.880 2.270 7.100 2.550 ;
        RECT  6.880 0.700 7.100 0.980 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.240 5.100 1.800 ;
        RECT  4.640 1.340 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.260 -0.280 5.540 0.760 ;
        RECT  6.300 -0.280 6.580 0.760 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.420 2.270 3.480 ;
        RECT  2.660 2.420 2.940 3.480 ;
        RECT  4.660 2.680 4.940 3.480 ;
        RECT  6.300 2.620 6.580 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.320 2.300 5.480 2.640 ;
        RECT  5.320 2.300 6.680 2.460 ;
        RECT  6.520 0.980 6.680 2.460 ;
        RECT  5.840 0.980 6.680 1.140 ;
        RECT  5.840 0.540 6.000 1.140 ;
        RECT  3.100 2.420 4.390 2.580 ;
        RECT  5.000 1.960 5.160 2.520 ;
        RECT  4.230 2.360 5.160 2.520 ;
        RECT  3.100 2.100 3.260 2.580 ;
        RECT  0.940 2.100 3.260 2.260 ;
        RECT  5.000 1.960 6.140 2.120 ;
        RECT  5.980 1.450 6.140 2.120 ;
        RECT  1.720 0.760 1.880 2.260 ;
        RECT  1.660 0.760 1.940 0.920 ;
        RECT  3.500 1.980 3.780 2.260 ;
        RECT  3.500 1.980 4.380 2.140 ;
        RECT  4.220 0.760 4.380 2.140 ;
        RECT  5.450 0.920 5.610 1.570 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  4.220 0.760 4.500 1.080 ;
        RECT  2.720 0.920 3.920 1.080 ;
        RECT  3.760 0.440 3.920 1.080 ;
        RECT  2.720 0.660 2.880 1.080 ;
        RECT  4.740 0.440 5.020 0.760 ;
        RECT  3.760 0.440 5.020 0.600 ;
        RECT  0.100 0.920 1.360 1.080 ;
        RECT  1.200 0.440 1.360 1.080 ;
        RECT  0.160 0.660 0.320 1.080 ;
        RECT  2.180 0.440 2.460 0.760 ;
        RECT  1.200 0.440 2.460 0.600 ;
    END
END OAI2222CHD

MACRO OAI2222EHD
    CLASS CORE ;
    FOREIGN OAI2222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.700 7.100 2.550 ;
        RECT  6.880 2.270 7.100 2.550 ;
        RECT  6.860 0.700 7.100 0.980 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.240 5.100 1.800 ;
        RECT  4.640 1.340 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.220 -0.280 5.500 0.760 ;
        RECT  6.280 -0.280 6.560 0.760 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.420 2.270 3.480 ;
        RECT  2.660 2.420 2.940 3.480 ;
        RECT  4.660 2.680 4.940 3.480 ;
        RECT  6.300 2.620 6.580 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.320 2.300 5.480 2.640 ;
        RECT  5.320 2.300 6.680 2.460 ;
        RECT  6.520 0.980 6.680 2.460 ;
        RECT  5.800 0.980 6.680 1.140 ;
        RECT  5.800 0.540 5.960 1.140 ;
        RECT  3.100 2.420 4.390 2.580 ;
        RECT  5.000 1.960 5.160 2.520 ;
        RECT  4.230 2.360 5.160 2.520 ;
        RECT  3.100 2.100 3.260 2.580 ;
        RECT  0.940 2.100 3.260 2.260 ;
        RECT  5.000 1.960 6.140 2.120 ;
        RECT  5.980 1.450 6.140 2.120 ;
        RECT  1.720 0.920 1.880 2.260 ;
        RECT  1.660 0.920 1.940 1.080 ;
        RECT  3.500 1.980 3.780 2.260 ;
        RECT  3.500 1.980 4.380 2.140 ;
        RECT  4.220 0.920 4.380 2.140 ;
        RECT  5.450 0.920 5.610 1.570 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  2.620 0.920 3.980 1.080 ;
        RECT  3.820 0.600 3.980 1.080 ;
        RECT  3.820 0.600 5.020 0.760 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OAI2222EHD

MACRO OAI2222HHD
    CLASS CORE ;
    FOREIGN OAI2222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.700 7.100 2.280 ;
        RECT  6.620 2.070 7.100 2.280 ;
        RECT  6.840 0.700 7.100 0.980 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.240 5.100 1.800 ;
        RECT  4.640 1.340 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.220 -0.280 5.500 0.760 ;
        RECT  6.260 -0.280 6.540 0.760 ;
        RECT  7.400 -0.280 7.680 0.760 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.420 2.270 3.480 ;
        RECT  2.660 2.420 2.940 3.480 ;
        RECT  4.550 2.680 4.830 3.480 ;
        RECT  6.100 2.620 6.380 3.480 ;
        RECT  7.170 2.430 7.450 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.320 2.300 5.540 2.760 ;
        RECT  5.320 2.300 6.460 2.460 ;
        RECT  6.300 1.750 6.460 2.460 ;
        RECT  6.460 0.980 6.620 1.910 ;
        RECT  5.800 0.980 6.620 1.140 ;
        RECT  5.800 0.540 5.960 1.140 ;
        RECT  3.100 2.420 4.390 2.580 ;
        RECT  5.000 1.960 5.160 2.520 ;
        RECT  4.230 2.360 5.160 2.520 ;
        RECT  3.100 2.100 3.260 2.580 ;
        RECT  0.940 2.100 3.260 2.260 ;
        RECT  5.000 1.960 6.140 2.120 ;
        RECT  5.980 1.450 6.140 2.120 ;
        RECT  1.720 0.920 1.880 2.260 ;
        RECT  1.660 0.920 1.940 1.080 ;
        RECT  3.500 1.980 3.780 2.260 ;
        RECT  3.500 1.980 4.380 2.140 ;
        RECT  4.220 0.920 4.380 2.140 ;
        RECT  5.450 0.920 5.610 1.570 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  2.620 0.920 3.980 1.080 ;
        RECT  3.820 0.600 3.980 1.080 ;
        RECT  3.820 0.600 5.020 0.760 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OAI2222HHD

MACRO OAI2222KHD
    CLASS CORE ;
    FOREIGN OAI2222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.620 2.100 8.000 2.300 ;
        RECT  6.780 0.740 8.160 0.940 ;
        RECT  7.300 0.740 7.500 2.300 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN D2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        END
    END D2
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.760 ;
        END
    END D1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 4.060 1.620 ;
        RECT  3.700 1.240 3.900 1.760 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.900 1.240 5.100 1.800 ;
        RECT  4.640 1.340 5.100 1.620 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.180 -0.280 3.460 0.760 ;
        RECT  5.220 -0.280 5.500 0.760 ;
        RECT  6.260 -0.280 6.540 0.760 ;
        RECT  7.300 -0.280 7.580 0.580 ;
        RECT  8.400 -0.280 8.680 0.580 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.420 2.270 3.480 ;
        RECT  2.660 2.420 2.940 3.480 ;
        RECT  4.690 2.580 4.970 3.480 ;
        RECT  6.100 2.620 6.380 3.480 ;
        RECT  7.170 2.620 7.450 3.480 ;
        RECT  8.270 2.620 8.550 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.320 2.300 5.480 2.760 ;
        RECT  5.320 2.300 6.460 2.460 ;
        RECT  6.300 1.750 6.460 2.460 ;
        RECT  6.460 0.980 6.620 1.910 ;
        RECT  5.800 0.980 6.620 1.140 ;
        RECT  5.800 0.540 5.960 1.140 ;
        RECT  3.100 2.420 4.390 2.580 ;
        RECT  5.000 1.960 5.160 2.420 ;
        RECT  4.230 2.260 5.160 2.420 ;
        RECT  3.100 2.100 3.260 2.580 ;
        RECT  0.940 2.100 3.260 2.260 ;
        RECT  5.000 1.960 6.140 2.120 ;
        RECT  5.980 1.450 6.140 2.120 ;
        RECT  1.720 0.920 1.880 2.260 ;
        RECT  1.660 0.920 1.940 1.080 ;
        RECT  3.500 1.940 3.780 2.260 ;
        RECT  3.500 1.940 4.380 2.100 ;
        RECT  4.220 0.920 4.380 2.100 ;
        RECT  5.450 0.920 5.610 1.570 ;
        RECT  4.220 0.920 5.610 1.080 ;
        RECT  2.620 0.920 3.980 1.080 ;
        RECT  3.820 0.600 3.980 1.080 ;
        RECT  3.820 0.600 5.020 0.760 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OAI2222KHD

MACRO OAI222BHD
    CLASS CORE ;
    FOREIGN OAI222BHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.870 4.300 2.280 ;
        RECT  1.880 2.120 4.300 2.280 ;
        RECT  3.460 0.870 4.300 1.030 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 1.340 3.910 1.620 ;
        RECT  3.700 1.240 3.900 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.800 ;
        RECT  3.260 1.340 3.500 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.210 1.900 1.800 ;
        RECT  1.650 1.390 1.900 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.730 1.390 1.100 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 -0.280 1.740 0.710 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.100 -0.280 0.380 1.000 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.980 2.620 3.260 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.280 2.440 0.560 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.940 0.550 4.300 0.710 ;
        RECT  0.900 0.870 2.780 1.030 ;
    END
END OAI222BHD

MACRO OAI222EHD
    CLASS CORE ;
    FOREIGN OAI222EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.880 5.500 2.340 ;
        RECT  5.280 2.060 5.500 2.340 ;
        RECT  5.280 0.880 5.500 1.160 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.710 ;
        RECT  4.700 -0.280 4.980 1.060 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.710 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.580 2.840 3.480 ;
        RECT  4.700 2.620 4.980 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.100 2.480 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.170 2.160 4.400 2.440 ;
        RECT  4.240 0.880 4.400 2.440 ;
        RECT  4.240 1.400 5.140 1.600 ;
        RECT  1.480 2.260 3.880 2.420 ;
        RECT  3.720 1.470 3.880 2.420 ;
        RECT  3.720 1.470 4.060 1.630 ;
        RECT  3.900 0.870 4.060 1.630 ;
        RECT  3.140 0.870 4.060 1.030 ;
        RECT  1.620 0.550 3.980 0.710 ;
        RECT  0.580 0.870 2.420 1.030 ;
    END
END OAI222EHD

MACRO OAI222HHD
    CLASS CORE ;
    FOREIGN OAI222HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.900 5.900 2.300 ;
        RECT  5.480 2.100 5.900 2.300 ;
        RECT  5.480 0.900 5.900 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.710 ;
        RECT  4.920 -0.280 5.200 0.860 ;
        RECT  6.000 -0.280 6.280 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.710 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.440 2.840 3.480 ;
        RECT  4.910 2.620 5.190 3.480 ;
        RECT  6.020 2.620 6.300 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.100 2.300 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.450 0.880 4.610 2.460 ;
        RECT  4.450 1.400 5.540 1.600 ;
        RECT  1.480 2.080 3.880 2.240 ;
        RECT  3.720 1.470 3.880 2.240 ;
        RECT  3.720 1.470 4.060 1.630 ;
        RECT  3.900 0.870 4.060 1.630 ;
        RECT  3.140 0.870 4.060 1.030 ;
        RECT  1.620 0.550 3.980 0.710 ;
        RECT  0.580 0.870 2.420 1.030 ;
    END
END OAI222HHD

MACRO OAI222KHD
    CLASS CORE ;
    FOREIGN OAI222KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.640 0.900 6.980 1.100 ;
        RECT  5.640 2.100 6.980 2.300 ;
        RECT  6.500 0.900 6.700 2.300 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.240 2.700 1.800 ;
        RECT  2.340 1.340 2.700 1.620 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.800 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.340 3.540 1.620 ;
        RECT  3.300 1.240 3.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.240 3.100 1.800 ;
        RECT  2.860 1.340 3.100 1.620 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.210 1.500 1.800 ;
        RECT  1.250 1.390 1.500 1.670 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.240 0.700 1.800 ;
        RECT  0.410 1.390 0.700 1.670 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.710 ;
        RECT  5.120 -0.280 5.400 0.580 ;
        RECT  6.160 -0.280 6.440 0.580 ;
        RECT  7.220 -0.280 7.500 0.580 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.710 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 2.490 2.840 3.480 ;
        RECT  5.120 2.620 5.400 3.480 ;
        RECT  6.180 2.620 6.460 3.480 ;
        RECT  7.220 2.620 7.500 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.100 2.350 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.660 0.880 4.820 2.380 ;
        RECT  4.660 1.400 5.960 1.600 ;
        RECT  4.620 0.880 4.820 1.160 ;
        RECT  1.480 2.080 4.060 2.240 ;
        RECT  3.900 0.870 4.060 2.240 ;
        RECT  3.140 0.870 4.060 1.030 ;
        RECT  1.620 0.550 3.980 0.710 ;
        RECT  0.580 0.870 2.420 1.030 ;
    END
END OAI222KHD

MACRO OAI22CHD
    CLASS CORE ;
    FOREIGN OAI22CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.940 2.100 1.900 2.300 ;
        RECT  1.700 0.950 1.900 2.300 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.620 -0.280 0.900 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.990 2.440 2.270 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 2.620 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 0.920 1.420 1.080 ;
        RECT  1.260 0.600 1.420 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.260 0.600 2.460 0.760 ;
    END
END OAI22CHD

MACRO OAI22EHD
    CLASS CORE ;
    FOREIGN OAI22EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.880 4.300 2.340 ;
        RECT  4.080 2.060 4.300 2.340 ;
        RECT  4.060 0.880 4.300 1.160 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.340 1.580 1.620 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.480 -0.280 3.760 1.060 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.020 2.420 2.300 3.480 ;
        RECT  3.500 2.620 3.780 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.970 2.160 3.160 2.440 ;
        RECT  3.000 0.880 3.160 2.440 ;
        RECT  3.000 1.420 3.940 1.580 ;
        RECT  1.020 2.100 2.780 2.260 ;
        RECT  2.620 0.920 2.780 2.260 ;
        RECT  1.700 0.920 2.780 1.080 ;
        RECT  0.100 0.920 1.500 1.080 ;
        RECT  1.340 0.600 1.500 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.340 0.600 2.580 0.760 ;
    END
END OAI22EHD

MACRO OAI22HHD
    CLASS CORE ;
    FOREIGN OAI22HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.900 4.300 2.300 ;
        RECT  3.880 2.100 4.300 2.300 ;
        RECT  3.880 0.900 4.300 1.100 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.340 1.580 1.620 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.320 -0.280 3.600 0.860 ;
        RECT  4.400 -0.280 4.680 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.020 2.420 2.300 3.480 ;
        RECT  3.310 2.620 3.590 3.480 ;
        RECT  4.420 2.620 4.700 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.850 0.840 3.010 2.460 ;
        RECT  2.850 1.420 3.940 1.580 ;
        RECT  1.020 2.100 2.620 2.260 ;
        RECT  2.460 0.920 2.620 2.260 ;
        RECT  1.700 0.920 2.620 1.080 ;
        RECT  0.100 0.920 1.500 1.080 ;
        RECT  1.340 0.600 1.500 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.340 0.600 2.580 0.760 ;
    END
END OAI22HHD

MACRO OAI22KHD
    CLASS CORE ;
    FOREIGN OAI22KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.040 0.900 5.380 1.100 ;
        RECT  4.040 2.100 5.380 2.300 ;
        RECT  4.900 0.900 5.100 2.300 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.800 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.800 ;
        RECT  0.860 1.340 1.100 1.620 ;
        END
    END B1
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.340 1.580 1.620 ;
        RECT  1.300 1.240 1.500 1.800 ;
        END
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.240 2.300 1.800 ;
        RECT  1.980 1.340 2.300 1.620 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.520 -0.280 3.800 0.580 ;
        RECT  4.560 -0.280 4.840 0.580 ;
        RECT  5.620 -0.280 5.900 0.580 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.020 2.420 2.300 3.480 ;
        RECT  3.520 2.620 3.800 3.480 ;
        RECT  4.580 2.620 4.860 3.480 ;
        RECT  5.620 2.620 5.900 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.100 2.420 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.050 2.060 3.280 2.340 ;
        RECT  3.050 0.880 3.210 2.340 ;
        RECT  3.050 1.420 4.360 1.580 ;
        RECT  3.020 0.880 3.210 1.160 ;
        RECT  1.020 2.100 2.620 2.260 ;
        RECT  2.460 0.920 2.620 2.260 ;
        RECT  1.700 0.920 2.620 1.080 ;
        RECT  0.100 0.920 1.500 1.080 ;
        RECT  1.340 0.600 1.500 1.080 ;
        RECT  0.100 0.860 0.380 1.080 ;
        RECT  1.340 0.600 2.580 0.760 ;
    END
END OAI22KHD

MACRO OR2B1CHD
    CLASS CORE ;
    FOREIGN OR2B1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.660 1.900 2.440 ;
        RECT  1.140 2.240 1.900 2.440 ;
        RECT  1.680 0.660 1.900 0.940 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.390 0.320 1.670 ;
        RECT  0.100 1.240 0.300 1.750 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.100 1.750 ;
        RECT  0.860 1.240 1.100 1.520 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.680 -0.280 0.960 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  0.680 2.800 1.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.280 0.980 2.440 ;
        RECT  0.820 1.920 0.980 2.440 ;
        RECT  0.100 2.220 0.380 2.440 ;
        RECT  0.820 1.920 1.540 2.080 ;
        RECT  1.320 1.480 1.540 2.080 ;
        RECT  1.360 0.800 1.520 2.080 ;
        RECT  0.100 0.800 1.520 0.960 ;
    END
END OR2B1CHD

MACRO OR2B1EHD
    CLASS CORE ;
    FOREIGN OR2B1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.710 2.700 2.480 ;
        RECT  2.480 2.200 2.700 2.480 ;
        RECT  2.480 0.710 2.700 0.990 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.140 1.540 1.420 ;
        RECT  1.300 1.140 1.500 1.650 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.450 0.300 1.960 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.800 -0.280 2.080 0.640 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.680 -0.280 0.840 0.720 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.960 2.520 2.120 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.680 2.440 0.840 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.920 1.920 2.260 2.080 ;
        RECT  2.100 0.820 2.260 2.080 ;
        RECT  2.100 1.390 2.340 1.670 ;
        RECT  1.140 0.820 2.260 0.980 ;
        RECT  0.160 2.120 0.380 2.720 ;
        RECT  0.160 2.120 0.680 2.280 ;
        RECT  0.520 0.880 0.680 2.280 ;
        RECT  0.520 1.390 1.000 1.670 ;
        RECT  0.160 0.880 0.680 1.040 ;
        RECT  0.160 0.440 0.380 1.040 ;
    END
END OR2B1EHD

MACRO OR2B1HHD
    CLASS CORE ;
    FOREIGN OR2B1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.850 0.770 3.150 2.350 ;
        RECT  2.700 2.050 3.150 2.350 ;
        RECT  2.670 0.770 3.150 1.070 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.140 1.540 1.420 ;
        RECT  1.300 1.140 1.500 1.650 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.450 0.300 1.960 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.800 -0.280 2.080 0.640 ;
        RECT  3.220 -0.280 3.500 0.580 ;
        RECT  0.000 -0.280 3.600 0.280 ;
        RECT  0.680 -0.280 0.840 0.720 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.180 2.520 2.340 3.480 ;
        RECT  3.280 2.480 3.440 3.480 ;
        RECT  0.000 2.920 3.600 3.480 ;
        RECT  0.160 2.350 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.140 1.920 2.480 2.080 ;
        RECT  2.320 0.820 2.480 2.080 ;
        RECT  2.320 1.390 2.560 1.670 ;
        RECT  1.140 0.820 2.480 0.980 ;
        RECT  0.680 2.310 0.900 2.630 ;
        RECT  0.680 1.390 0.840 2.630 ;
        RECT  0.520 1.390 1.000 1.670 ;
        RECT  0.520 0.880 0.680 1.670 ;
        RECT  0.160 0.880 0.680 1.040 ;
        RECT  0.160 0.440 0.380 1.040 ;
    END
END OR2B1HHD

MACRO OR2B1KHD
    CLASS CORE ;
    FOREIGN OR2B1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.490 0.800 5.250 1.300 ;
        RECT  4.670 0.780 4.830 1.300 ;
        RECT  4.750 0.800 5.250 2.400 ;
        RECT  3.660 1.900 5.250 2.400 ;
        RECT  3.550 0.780 3.710 1.300 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.050 1.520 2.330 1.680 ;
        RECT  2.100 1.520 2.300 2.050 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.450 0.300 1.960 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.800 -0.280 2.080 0.640 ;
        RECT  2.960 -0.280 3.240 0.640 ;
        RECT  4.020 -0.280 4.300 0.640 ;
        RECT  5.220 -0.280 5.500 0.640 ;
        RECT  0.000 -0.280 5.600 0.280 ;
        RECT  0.680 -0.280 0.840 0.720 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.960 2.560 2.240 3.480 ;
        RECT  3.140 2.560 3.420 3.480 ;
        RECT  4.180 2.560 4.460 3.480 ;
        RECT  5.220 2.560 5.500 3.480 ;
        RECT  0.000 2.920 5.600 3.480 ;
        RECT  0.160 2.330 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.120 2.240 3.020 2.400 ;
        RECT  2.860 1.720 3.020 2.400 ;
        RECT  2.860 1.720 3.280 1.880 ;
        RECT  3.120 0.820 3.280 1.880 ;
        RECT  1.140 0.820 3.280 0.980 ;
        RECT  0.680 2.330 0.900 2.610 ;
        RECT  0.680 1.140 0.840 2.610 ;
        RECT  0.680 1.200 2.860 1.360 ;
        RECT  0.520 0.880 0.680 1.300 ;
        RECT  0.160 0.880 0.680 1.040 ;
        RECT  0.160 0.440 0.380 1.040 ;
    END
END OR2B1KHD

MACRO OR2CHD
    CLASS CORE ;
    FOREIGN OR2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.650 1.900 2.500 ;
        RECT  1.680 2.220 1.900 2.500 ;
        RECT  1.680 0.650 1.900 0.930 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.130 0.320 1.410 ;
        RECT  0.100 1.130 0.300 1.670 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 1.960 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.060 -0.280 1.340 0.400 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  1.020 2.440 1.300 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.120 0.380 2.340 ;
        RECT  0.100 2.120 1.520 2.280 ;
        RECT  1.360 0.810 1.520 2.280 ;
        RECT  0.560 0.810 1.520 0.970 ;
    END
END OR2CHD

MACRO OR2EHD
    CLASS CORE ;
    FOREIGN OR2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.650 1.900 2.500 ;
        RECT  1.680 2.220 1.900 2.500 ;
        RECT  1.680 0.650 1.900 0.930 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.140 0.320 1.420 ;
        RECT  0.100 1.130 0.300 1.670 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.420 1.100 1.960 ;
        RECT  0.880 1.520 1.100 1.800 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.060 -0.280 1.340 0.400 ;
        RECT  0.000 -0.280 2.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.000 3.480 ;
        RECT  1.100 2.620 1.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.120 0.380 2.340 ;
        RECT  0.100 2.120 1.520 2.280 ;
        RECT  1.360 0.800 1.520 2.280 ;
        RECT  0.560 0.800 1.520 0.960 ;
    END
END OR2EHD

MACRO OR2HHD
    CLASS CORE ;
    FOREIGN OR2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 0.650 2.300 2.500 ;
        RECT  1.960 2.220 2.300 2.500 ;
        RECT  1.960 0.650 2.300 0.930 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.300 0.320 1.580 ;
        RECT  0.100 1.130 0.300 1.670 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.130 1.100 1.670 ;
        RECT  0.940 1.100 1.100 1.670 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  2.480 -0.280 2.700 0.640 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.480 2.560 2.700 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.380 2.620 1.660 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.500 2.120 1.800 2.280 ;
        RECT  1.640 0.600 1.800 2.280 ;
        RECT  0.780 0.600 1.800 0.760 ;
    END
END OR2HHD

MACRO OR2KHD
    CLASS CORE ;
    FOREIGN OR2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.740 3.100 2.360 ;
        RECT  2.880 2.080 3.100 2.360 ;
        RECT  3.920 0.740 4.300 1.020 ;
        RECT  2.900 1.240 4.300 1.560 ;
        RECT  4.100 0.740 4.300 2.360 ;
        RECT  3.920 2.080 4.300 2.360 ;
        RECT  2.880 0.740 3.100 1.020 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.080 1.500 1.600 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.080 1.460 2.280 1.740 ;
        RECT  2.120 1.460 2.280 2.280 ;
        RECT  0.500 2.120 2.280 2.280 ;
        RECT  0.500 1.460 0.700 2.420 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.260 -0.280 1.540 0.580 ;
        RECT  2.300 -0.280 2.580 0.580 ;
        RECT  3.340 -0.280 3.620 0.580 ;
        RECT  4.380 -0.280 4.660 0.580 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.760 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 2.800 2.480 3.480 ;
        RECT  3.340 2.620 3.620 3.480 ;
        RECT  4.380 2.620 4.660 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.180 2.580 0.460 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.260 2.480 2.720 2.640 ;
        RECT  2.560 0.760 2.720 2.640 ;
        RECT  0.660 0.760 2.720 0.920 ;
        RECT  1.840 0.520 2.000 0.920 ;
        RECT  0.660 0.700 0.940 0.920 ;
    END
END OR2KHD

MACRO OR3B1CHD
    CLASS CORE ;
    FOREIGN OR3B1CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.600 3.100 2.420 ;
        RECT  2.880 2.140 3.100 2.420 ;
        RECT  2.880 0.600 3.100 0.880 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.140 1.900 1.650 ;
        RECT  1.580 1.140 1.900 1.420 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.460 2.300 1.960 ;
        RECT  2.060 1.460 2.300 1.740 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.550 0.300 2.060 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.400 ;
        RECT  2.360 -0.280 2.520 0.640 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.160 -0.280 0.320 1.240 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.300 2.460 2.580 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.160 2.340 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.080 2.120 2.660 2.280 ;
        RECT  2.500 0.820 2.660 2.280 ;
        RECT  1.080 1.840 1.300 2.280 ;
        RECT  2.500 1.390 2.740 1.670 ;
        RECT  1.320 0.820 2.660 0.980 ;
        RECT  1.320 0.560 1.480 0.980 ;
        RECT  0.610 0.560 1.480 0.720 ;
        RECT  0.610 0.440 0.890 0.720 ;
        RECT  0.680 0.960 0.840 2.620 ;
        RECT  0.680 1.390 1.030 1.670 ;
    END
END OR3B1CHD

MACRO OR3B1EHD
    CLASS CORE ;
    FOREIGN OR3B1EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 0.600 3.100 2.420 ;
        RECT  2.880 2.140 3.100 2.420 ;
        RECT  2.880 0.600 3.100 0.880 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.140 1.900 1.650 ;
        RECT  1.580 1.140 1.900 1.420 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.460 2.300 1.960 ;
        RECT  2.060 1.460 2.300 1.740 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.550 0.300 2.060 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.220 -0.280 1.500 0.400 ;
        RECT  2.360 -0.280 2.520 0.640 ;
        RECT  0.000 -0.280 3.200 0.280 ;
        RECT  0.160 -0.280 0.320 1.240 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.360 2.460 2.520 3.480 ;
        RECT  0.000 2.920 3.200 3.480 ;
        RECT  0.160 2.320 0.320 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.080 2.120 2.660 2.280 ;
        RECT  2.500 0.820 2.660 2.280 ;
        RECT  1.080 1.840 1.270 2.280 ;
        RECT  2.500 1.390 2.740 1.670 ;
        RECT  1.320 0.820 2.660 0.980 ;
        RECT  1.320 0.560 1.480 0.980 ;
        RECT  0.610 0.560 1.480 0.720 ;
        RECT  0.610 0.440 0.890 0.720 ;
        RECT  0.680 0.960 0.840 2.600 ;
        RECT  0.680 1.390 1.030 1.670 ;
    END
END OR3B1EHD

MACRO OR3B1HHD
    CLASS CORE ;
    FOREIGN OR3B1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.100 0.660 4.300 2.300 ;
        RECT  3.880 2.100 4.300 2.300 ;
        RECT  3.680 0.660 4.300 0.860 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.380 1.360 2.540 1.940 ;
        RECT  1.300 1.780 2.540 1.940 ;
        RECT  2.550 1.060 2.770 1.520 ;
        RECT  2.380 1.360 2.770 1.520 ;
        RECT  1.300 1.460 1.590 1.940 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 2.120 2.880 2.280 ;
        RECT  2.720 1.960 3.240 2.120 ;
        RECT  3.080 1.460 3.240 2.120 ;
        RECT  0.900 1.460 1.100 2.280 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.550 0.300 2.060 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.740 -0.280 2.020 0.580 ;
        RECT  2.920 -0.280 3.200 0.580 ;
        RECT  4.360 -0.280 4.640 0.400 ;
        RECT  0.000 -0.280 4.800 0.280 ;
        RECT  0.680 -0.280 0.840 0.880 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.360 2.620 3.640 3.480 ;
        RECT  4.400 2.620 4.680 3.480 ;
        RECT  0.000 2.920 4.800 3.480 ;
        RECT  0.680 2.620 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.020 2.600 3.200 2.760 ;
        RECT  3.040 2.280 3.200 2.760 ;
        RECT  3.040 2.280 3.720 2.440 ;
        RECT  3.560 1.120 3.720 2.440 ;
        RECT  3.260 1.120 3.720 1.280 ;
        RECT  3.260 0.740 3.420 1.280 ;
        RECT  1.180 0.740 3.420 0.900 ;
        RECT  1.180 0.700 1.460 0.900 ;
        RECT  0.100 2.280 0.380 2.540 ;
        RECT  0.100 2.280 0.640 2.440 ;
        RECT  0.480 1.100 0.640 2.440 ;
        RECT  1.920 1.100 2.080 1.620 ;
        RECT  0.160 1.100 2.080 1.260 ;
        RECT  0.160 0.600 0.320 1.260 ;
    END
END OR3B1HHD

MACRO OR3B2CHD
    CLASS CORE ;
    FOREIGN OR3B2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.500 2.700 2.320 ;
        RECT  1.300 2.120 2.700 2.320 ;
        RECT  2.150 0.500 2.700 0.700 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.650 0.320 1.930 ;
        RECT  0.100 1.520 0.300 2.060 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.220 1.620 ;
        RECT  0.900 1.220 1.100 1.760 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.440 1.900 1.960 ;
        RECT  1.560 1.560 1.900 1.840 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.740 -0.280 0.900 0.640 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 2.520 2.140 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.840 2.280 1.000 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.100 2.380 0.640 2.540 ;
        RECT  0.480 0.900 0.640 2.540 ;
        RECT  2.170 0.900 2.330 1.620 ;
        RECT  0.100 0.900 0.640 1.140 ;
        RECT  0.100 0.900 2.330 1.060 ;
    END
END OR3B2CHD

MACRO OR3B2EHD
    CLASS CORE ;
    FOREIGN OR3B2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.600 3.900 2.420 ;
        RECT  3.680 2.140 3.900 2.420 ;
        RECT  3.680 0.600 3.900 0.880 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.460 3.100 1.960 ;
        RECT  2.860 1.460 3.100 1.740 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.600 0.320 1.880 ;
        RECT  0.100 1.600 0.300 2.110 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.160 1.740 ;
        RECT  0.900 1.400 1.100 1.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.620 0.940 0.900 1.100 ;
        RECT  2.020 -0.280 2.300 0.400 ;
        RECT  3.160 -0.280 3.320 0.640 ;
        RECT  0.000 -0.280 4.000 0.280 ;
        RECT  0.680 -0.280 0.840 1.100 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 2.560 3.380 3.480 ;
        RECT  0.000 2.920 4.000 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.730 2.600 2.910 2.760 ;
        RECT  2.750 2.220 2.910 2.760 ;
        RECT  2.750 2.220 3.460 2.380 ;
        RECT  3.300 0.820 3.460 2.380 ;
        RECT  3.300 1.390 3.540 1.670 ;
        RECT  2.120 0.820 3.460 0.980 ;
        RECT  2.120 0.560 2.280 0.980 ;
        RECT  1.410 0.560 2.280 0.720 ;
        RECT  1.410 0.440 1.690 0.720 ;
        RECT  0.100 2.280 0.380 2.540 ;
        RECT  0.100 2.280 2.540 2.440 ;
        RECT  2.380 1.140 2.540 2.440 ;
        RECT  0.520 1.280 0.680 2.440 ;
        RECT  0.160 1.280 0.680 1.440 ;
        RECT  2.320 1.140 2.540 1.420 ;
        RECT  0.160 0.880 0.380 1.440 ;
        RECT  1.280 1.960 1.560 2.120 ;
        RECT  1.380 0.960 1.540 2.120 ;
        RECT  1.380 1.460 1.830 1.740 ;
        RECT  1.240 0.960 1.540 1.240 ;
    END
END OR3B2EHD

MACRO OR3B2HHD
    CLASS CORE ;
    FOREIGN OR3B2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.140 2.060 5.300 2.340 ;
        RECT  5.300 0.660 5.500 2.300 ;
        RECT  5.080 2.100 5.500 2.300 ;
        RECT  4.880 0.660 5.500 0.860 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.520 2.340 1.680 ;
        RECT  2.100 2.120 4.080 2.280 ;
        RECT  3.920 1.960 4.440 2.120 ;
        RECT  4.280 1.460 4.440 2.120 ;
        RECT  2.100 1.520 2.300 2.280 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.550 0.300 2.060 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.160 1.740 ;
        RECT  0.900 1.400 1.100 1.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.820 -0.280 2.100 0.400 ;
        RECT  2.940 -0.280 3.220 0.400 ;
        RECT  4.320 -0.280 4.600 0.420 ;
        RECT  5.560 -0.280 5.840 0.400 ;
        RECT  0.000 -0.280 6.000 0.280 ;
        RECT  0.680 -0.280 0.840 0.880 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.800 2.800 2.080 3.480 ;
        RECT  4.560 2.620 4.840 3.480 ;
        RECT  5.600 2.620 5.880 3.480 ;
        RECT  0.000 2.920 6.000 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.220 2.600 4.400 2.760 ;
        RECT  4.240 2.280 4.400 2.760 ;
        RECT  4.240 2.280 4.920 2.440 ;
        RECT  4.760 1.120 4.920 2.440 ;
        RECT  4.460 1.120 4.920 1.280 ;
        RECT  4.460 0.740 4.620 1.280 ;
        RECT  3.440 0.740 4.620 0.900 ;
        RECT  3.440 0.560 3.600 0.900 ;
        RECT  2.380 0.560 3.600 0.720 ;
        RECT  2.380 0.440 2.660 0.720 ;
        RECT  0.100 2.380 1.880 2.540 ;
        RECT  1.720 1.200 1.880 2.540 ;
        RECT  0.100 2.300 0.680 2.540 ;
        RECT  0.520 1.080 0.680 2.540 ;
        RECT  2.620 1.780 3.740 1.940 ;
        RECT  3.580 1.360 3.740 1.940 ;
        RECT  2.620 1.200 2.780 1.940 ;
        RECT  3.580 1.360 3.970 1.520 ;
        RECT  3.750 1.060 3.970 1.520 ;
        RECT  1.720 1.200 2.780 1.360 ;
        RECT  0.160 1.080 0.680 1.240 ;
        RECT  0.160 0.600 0.320 1.240 ;
        RECT  1.280 2.060 1.560 2.220 ;
        RECT  1.380 0.880 1.540 2.220 ;
        RECT  3.120 0.880 3.280 1.620 ;
        RECT  1.270 0.880 3.280 1.040 ;
        RECT  1.270 0.600 1.430 1.040 ;
    END
END OR3B2HHD

MACRO OR3B2KHD
    CLASS CORE ;
    FOREIGN OR3B2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.980 2.100 5.180 2.760 ;
        RECT  4.860 2.600 5.180 2.760 ;
        RECT  5.020 0.660 5.220 1.100 ;
        RECT  5.020 0.900 6.300 1.100 ;
        RECT  5.960 2.020 6.300 2.300 ;
        RECT  6.100 0.900 6.300 2.300 ;
        RECT  4.980 2.100 6.300 2.300 ;
        RECT  4.800 0.660 5.220 0.860 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.520 2.300 2.280 ;
        RECT  3.700 1.910 3.860 2.280 ;
        RECT  2.100 2.120 3.860 2.280 ;
        RECT  4.200 1.460 4.360 2.070 ;
        RECT  3.700 1.910 4.360 2.070 ;
        RECT  1.980 1.520 2.300 1.740 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.550 0.320 1.830 ;
        RECT  0.100 1.550 0.300 2.060 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.460 1.110 1.740 ;
        RECT  0.900 1.130 1.100 1.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.740 -0.280 2.020 0.400 ;
        RECT  2.860 -0.280 3.140 0.400 ;
        RECT  4.240 -0.280 4.520 0.420 ;
        RECT  5.420 -0.280 5.580 0.640 ;
        RECT  6.480 -0.280 6.640 0.680 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.680 -0.280 0.840 0.880 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.720 2.800 2.000 3.480 ;
        RECT  4.380 2.560 4.540 3.480 ;
        RECT  5.380 2.620 5.660 3.480 ;
        RECT  6.420 2.620 6.700 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.140 2.600 4.180 2.760 ;
        RECT  4.020 2.230 4.180 2.760 ;
        RECT  4.020 2.230 4.820 2.390 ;
        RECT  4.660 1.120 4.820 2.390 ;
        RECT  4.660 1.390 4.840 1.670 ;
        RECT  4.380 1.120 4.820 1.280 ;
        RECT  4.380 0.740 4.540 1.280 ;
        RECT  3.360 0.740 4.540 0.900 ;
        RECT  3.360 0.560 3.520 0.900 ;
        RECT  2.300 0.560 3.520 0.720 ;
        RECT  2.300 0.440 2.580 0.720 ;
        RECT  0.100 2.440 1.820 2.600 ;
        RECT  1.660 1.200 1.820 2.600 ;
        RECT  0.100 2.380 0.680 2.600 ;
        RECT  0.520 1.080 0.680 2.600 ;
        RECT  2.540 1.780 3.520 1.940 ;
        RECT  3.360 1.360 3.520 1.940 ;
        RECT  2.540 1.200 2.700 1.940 ;
        RECT  3.360 1.360 3.890 1.520 ;
        RECT  3.670 1.060 3.890 1.520 ;
        RECT  1.660 1.200 2.700 1.360 ;
        RECT  0.160 1.080 0.680 1.240 ;
        RECT  0.160 0.600 0.320 1.240 ;
        RECT  1.270 2.000 1.460 2.280 ;
        RECT  1.270 0.600 1.430 2.280 ;
        RECT  3.040 0.880 3.200 1.620 ;
        RECT  1.270 0.880 3.200 1.040 ;
    END
END OR3B2KHD

MACRO OR3CHD
    CLASS CORE ;
    FOREIGN OR3CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.720 2.700 2.500 ;
        RECT  2.480 2.220 2.700 2.500 ;
        RECT  2.480 0.720 2.700 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.120 1.100 1.640 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.420 1.900 1.960 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.820 2.620 2.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.660 2.300 2.320 2.460 ;
        RECT  2.160 0.660 2.320 2.460 ;
        RECT  2.160 1.220 2.340 1.500 ;
        RECT  0.100 0.660 2.320 0.820 ;
    END
END OR3CHD

MACRO OR3EHD
    CLASS CORE ;
    FOREIGN OR3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 0.720 2.700 2.500 ;
        RECT  2.480 2.220 2.700 2.500 ;
        RECT  2.480 0.720 2.700 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.120 1.120 1.400 ;
        RECT  0.900 1.120 1.100 1.640 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.420 1.900 1.960 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.420 0.700 1.960 ;
        RECT  0.480 1.460 0.700 1.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.860 -0.280 2.140 0.400 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  1.860 2.620 2.140 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.660 2.300 2.310 2.460 ;
        RECT  2.150 0.660 2.310 2.460 ;
        RECT  2.150 1.340 2.340 1.620 ;
        RECT  0.100 0.660 2.310 0.820 ;
    END
END OR3EHD

MACRO OR3HHD
    CLASS CORE ;
    FOREIGN OR3HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.700 0.720 3.900 2.500 ;
        RECT  3.560 2.220 3.900 2.500 ;
        RECT  3.560 0.720 3.900 1.000 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.040 0.900 2.300 1.100 ;
        RECT  2.100 0.900 2.300 1.560 ;
        RECT  1.040 0.900 1.260 1.340 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.740 1.460 2.900 2.280 ;
        RECT  0.500 2.120 2.900 2.280 ;
        RECT  0.500 1.420 0.700 2.360 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.420 1.900 1.960 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 -0.280 3.200 0.400 ;
        RECT  4.020 -0.280 4.300 0.580 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  1.740 -0.280 2.020 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 2.800 3.200 3.480 ;
        RECT  4.020 2.620 4.300 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.180 2.580 0.460 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.700 2.480 3.400 2.640 ;
        RECT  3.240 0.560 3.400 2.640 ;
        RECT  3.240 1.400 3.540 1.680 ;
        RECT  1.180 0.560 3.400 0.720 ;
    END
END OR3HHD

MACRO QDBAHEHD
    CLASS CORE ;
    FOREIGN QDBAHEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END GB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.850 5.510 1.130 ;
        RECT  5.300 1.840 5.510 2.120 ;
        RECT  5.300 0.850 5.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.980 ;
        RECT  5.890 -0.280 6.170 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.850 2.800 6.130 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 0.820 5.030 2.440 ;
        RECT  4.030 1.200 4.310 1.420 ;
        RECT  4.030 1.200 5.090 1.360 ;
        RECT  4.810 0.820 5.090 1.360 ;
        RECT  3.050 2.480 4.630 2.640 ;
        RECT  4.470 1.690 4.630 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.820 3.850 2.320 ;
        RECT  3.690 0.820 3.970 0.980 ;
        RECT  0.100 2.300 1.010 2.460 ;
        RECT  0.850 0.580 1.010 2.460 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.850 0.580 2.370 0.740 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  1.290 2.300 2.870 2.460 ;
        RECT  2.710 1.380 2.870 2.460 ;
        RECT  1.290 0.900 1.450 2.460 ;
        RECT  1.290 0.900 1.570 1.120 ;
        RECT  2.330 1.850 2.550 2.130 ;
        RECT  2.390 0.940 2.550 2.130 ;
        RECT  2.330 0.940 2.610 1.100 ;
    END
END QDBAHEHD

MACRO QDBAHHHD
    CLASS CORE ;
    FOREIGN QDBAHHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN GB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END GB
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.850 6.030 1.130 ;
        RECT  5.700 1.840 6.030 2.120 ;
        RECT  5.700 0.850 5.900 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.980 ;
        RECT  5.290 -0.280 5.570 0.580 ;
        RECT  6.330 -0.280 6.610 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.290 2.620 5.570 3.480 ;
        RECT  6.330 2.620 6.610 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 0.820 5.030 2.440 ;
        RECT  4.030 1.200 4.310 1.420 ;
        RECT  4.030 1.200 5.090 1.360 ;
        RECT  4.810 0.820 5.090 1.360 ;
        RECT  3.050 2.480 4.700 2.640 ;
        RECT  4.540 1.520 4.700 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.820 3.850 2.320 ;
        RECT  3.690 0.820 3.970 0.980 ;
        RECT  0.100 2.300 1.010 2.460 ;
        RECT  0.850 0.580 1.010 2.460 ;
        RECT  0.100 2.220 0.380 2.460 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.850 0.580 2.370 0.740 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  1.290 2.300 2.890 2.460 ;
        RECT  2.730 1.440 2.890 2.460 ;
        RECT  1.290 1.020 1.450 2.460 ;
        RECT  1.270 1.020 1.550 1.180 ;
        RECT  2.330 1.840 2.550 2.120 ;
        RECT  2.390 0.960 2.550 2.120 ;
    END
END QDBAHHHD

MACRO QDFFCHD
    CLASS CORE ;
    FOREIGN QDFFCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.780 ;
        RECT  1.180 1.310 1.500 1.590 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 0.440 7.900 2.120 ;
        RECT  7.680 1.840 7.900 2.120 ;
        RECT  7.620 0.440 7.900 0.660 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.280 -0.280 1.560 0.400 ;
        RECT  4.840 -0.280 5.120 0.420 ;
        RECT  6.320 -0.280 6.600 0.420 ;
        RECT  7.100 -0.280 7.380 0.600 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.800 1.660 3.480 ;
        RECT  4.710 2.800 4.990 3.480 ;
        RECT  5.760 2.800 6.500 3.480 ;
        RECT  7.100 2.060 7.460 2.280 ;
        RECT  7.220 2.060 7.460 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.720 2.540 7.060 2.760 ;
        RECT  2.800 2.600 3.790 2.760 ;
        RECT  3.630 2.160 3.790 2.760 ;
        RECT  5.850 2.480 6.880 2.640 ;
        RECT  2.800 0.460 2.960 2.760 ;
        RECT  6.720 0.920 6.880 2.760 ;
        RECT  5.850 1.860 6.010 2.640 ;
        RECT  2.380 2.300 2.960 2.460 ;
        RECT  3.630 2.160 4.170 2.320 ;
        RECT  4.010 1.860 4.170 2.320 ;
        RECT  4.010 1.860 6.010 2.020 ;
        RECT  6.710 0.920 7.040 1.140 ;
        RECT  2.680 0.460 2.960 0.680 ;
        RECT  6.260 0.580 6.420 2.120 ;
        RECT  6.260 1.340 6.560 1.620 ;
        RECT  5.720 0.580 6.420 0.740 ;
        RECT  3.120 2.180 3.470 2.440 ;
        RECT  3.120 0.460 3.280 2.440 ;
        RECT  5.920 1.140 6.080 1.660 ;
        RECT  3.760 1.140 6.080 1.300 ;
        RECT  3.760 0.460 3.920 1.300 ;
        RECT  3.120 0.460 3.920 0.620 ;
        RECT  5.280 0.580 5.560 0.980 ;
        RECT  4.080 0.580 5.560 0.740 ;
        RECT  4.080 0.460 4.680 0.740 ;
        RECT  4.040 2.480 4.570 2.640 ;
        RECT  5.280 2.180 5.560 2.520 ;
        RECT  4.410 2.360 5.560 2.520 ;
        RECT  3.440 1.460 3.840 1.980 ;
        RECT  3.440 1.460 5.420 1.620 ;
        RECT  3.440 0.840 3.600 1.980 ;
        RECT  0.600 1.700 0.760 2.210 ;
        RECT  2.480 0.880 2.640 2.080 ;
        RECT  0.580 0.440 0.740 1.860 ;
        RECT  2.360 0.440 2.520 1.040 ;
        RECT  0.580 0.560 1.880 0.720 ;
        RECT  1.720 0.440 2.520 0.600 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.000 0.840 2.160 2.320 ;
        RECT  2.000 1.380 2.300 1.660 ;
        RECT  0.900 2.400 1.820 2.560 ;
        RECT  1.660 0.920 1.820 2.560 ;
        RECT  0.900 0.920 1.820 1.080 ;
    END
END QDFFCHD

MACRO QDFFEHD
    CLASS CORE ;
    FOREIGN QDFFEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.780 ;
        RECT  1.170 1.350 1.500 1.630 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.440 7.500 2.120 ;
        RECT  7.160 1.840 7.500 2.120 ;
        RECT  7.100 0.440 7.500 0.660 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.190 -0.280 1.470 0.400 ;
        RECT  4.840 -0.280 5.120 0.420 ;
        RECT  6.320 -0.280 6.600 0.420 ;
        RECT  7.680 -0.280 7.900 0.660 ;
        RECT  0.000 -0.280 8.000 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.380 2.800 1.660 3.480 ;
        RECT  4.710 2.800 4.990 3.480 ;
        RECT  5.760 2.800 6.480 3.480 ;
        RECT  7.620 2.620 7.900 3.480 ;
        RECT  0.000 2.920 8.000 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.720 2.540 7.040 2.760 ;
        RECT  2.800 2.600 3.790 2.760 ;
        RECT  3.630 2.160 3.790 2.760 ;
        RECT  6.700 2.540 7.040 2.720 ;
        RECT  5.850 2.480 6.880 2.640 ;
        RECT  2.800 0.460 2.960 2.760 ;
        RECT  6.720 0.860 6.880 2.760 ;
        RECT  5.850 1.860 6.010 2.640 ;
        RECT  2.380 2.300 2.960 2.460 ;
        RECT  3.630 2.160 4.170 2.320 ;
        RECT  4.010 1.860 4.170 2.320 ;
        RECT  4.010 1.860 6.010 2.020 ;
        RECT  6.710 0.860 7.040 1.080 ;
        RECT  2.680 0.460 2.960 0.680 ;
        RECT  6.260 0.580 6.420 2.080 ;
        RECT  6.260 1.340 6.560 1.620 ;
        RECT  5.720 0.580 6.420 0.740 ;
        RECT  3.120 2.180 3.470 2.440 ;
        RECT  3.120 0.460 3.280 2.440 ;
        RECT  5.920 1.140 6.080 1.660 ;
        RECT  3.760 1.140 6.080 1.300 ;
        RECT  3.760 0.460 3.920 1.300 ;
        RECT  3.120 0.460 3.920 0.620 ;
        RECT  5.280 0.580 5.560 0.980 ;
        RECT  4.080 0.580 5.560 0.740 ;
        RECT  4.080 0.460 4.680 0.740 ;
        RECT  4.040 2.480 4.570 2.640 ;
        RECT  5.280 2.180 5.560 2.520 ;
        RECT  4.410 2.360 5.560 2.520 ;
        RECT  3.440 1.460 3.840 1.980 ;
        RECT  3.440 1.460 5.420 1.620 ;
        RECT  3.440 0.840 3.600 1.980 ;
        RECT  0.600 1.720 0.760 2.210 ;
        RECT  2.480 0.880 2.640 2.080 ;
        RECT  0.580 0.440 0.740 1.880 ;
        RECT  2.360 0.440 2.520 1.040 ;
        RECT  0.580 0.560 1.820 0.720 ;
        RECT  1.660 0.440 2.520 0.600 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.000 0.760 2.160 2.320 ;
        RECT  2.000 1.380 2.300 1.660 ;
        RECT  0.860 2.380 1.820 2.540 ;
        RECT  1.660 0.920 1.820 2.540 ;
        RECT  0.900 0.920 1.820 1.080 ;
    END
END QDFFEHD

MACRO QDFFHHD
    CLASS CORE ;
    FOREIGN QDFFHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.350 1.540 1.630 ;
        RECT  1.300 1.240 1.500 1.780 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.880 7.500 2.120 ;
        RECT  6.990 1.840 7.500 2.120 ;
        RECT  6.990 0.880 7.500 1.160 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.400 -0.280 1.680 0.400 ;
        RECT  5.050 -0.280 5.330 0.420 ;
        RECT  6.410 -0.280 6.690 0.580 ;
        RECT  7.450 -0.280 7.730 0.580 ;
        RECT  0.000 -0.280 8.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.590 2.800 1.870 3.480 ;
        RECT  4.840 2.800 5.120 3.480 ;
        RECT  6.410 2.620 6.690 3.480 ;
        RECT  7.450 2.620 7.730 3.480 ;
        RECT  0.000 2.920 8.400 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.010 2.600 4.000 2.760 ;
        RECT  3.840 2.160 4.000 2.760 ;
        RECT  3.010 0.460 3.170 2.760 ;
        RECT  5.970 2.300 8.190 2.460 ;
        RECT  8.030 0.910 8.190 2.460 ;
        RECT  2.590 2.300 3.170 2.460 ;
        RECT  5.570 2.220 6.130 2.380 ;
        RECT  3.840 2.160 4.380 2.320 ;
        RECT  5.570 2.030 5.730 2.380 ;
        RECT  4.220 2.030 5.730 2.190 ;
        RECT  2.890 0.460 3.170 0.680 ;
        RECT  5.890 1.840 6.420 2.060 ;
        RECT  6.260 1.000 6.420 2.060 ;
        RECT  6.260 1.340 6.830 1.620 ;
        RECT  6.050 1.000 6.420 1.160 ;
        RECT  6.050 0.440 6.210 1.160 ;
        RECT  5.850 0.440 6.210 0.600 ;
        RECT  3.330 2.180 3.680 2.440 ;
        RECT  3.330 0.460 3.490 2.440 ;
        RECT  5.840 1.350 6.060 1.630 ;
        RECT  3.970 1.350 6.060 1.510 ;
        RECT  3.970 0.460 4.130 1.510 ;
        RECT  3.330 0.460 4.130 0.620 ;
        RECT  4.730 0.940 5.810 1.100 ;
        RECT  4.730 0.460 4.890 1.100 ;
        RECT  4.290 0.460 4.890 0.740 ;
        RECT  5.250 2.540 5.810 2.700 ;
        RECT  4.250 2.480 4.780 2.640 ;
        RECT  5.250 2.360 5.410 2.700 ;
        RECT  4.620 2.360 5.410 2.520 ;
        RECT  3.650 1.680 4.050 1.980 ;
        RECT  3.650 1.680 5.630 1.840 ;
        RECT  3.650 0.840 3.810 1.980 ;
        RECT  0.600 0.560 0.760 2.170 ;
        RECT  2.690 0.880 2.850 2.080 ;
        RECT  2.570 0.440 2.730 1.040 ;
        RECT  0.600 0.560 2.030 0.720 ;
        RECT  1.870 0.440 2.730 0.600 ;
        RECT  2.210 0.760 2.370 2.320 ;
        RECT  2.210 1.380 2.510 1.660 ;
        RECT  1.110 2.150 2.030 2.310 ;
        RECT  1.870 0.920 2.030 2.310 ;
        RECT  1.110 0.920 2.030 1.080 ;
    END
END QDFFHHD

MACRO QDFFKHD
    CLASS CORE ;
    FOREIGN QDFFKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.240 1.900 1.780 ;
        RECT  1.660 1.350 1.900 1.630 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 0.880 8.500 1.160 ;
        RECT  7.300 1.840 8.500 2.120 ;
        RECT  7.700 0.880 7.900 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.280 2.120 0.400 ;
        RECT  5.300 -0.280 5.580 0.420 ;
        RECT  6.720 -0.280 7.000 0.580 ;
        RECT  7.760 -0.280 8.040 0.580 ;
        RECT  8.800 -0.280 9.080 0.580 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 2.800 2.120 3.480 ;
        RECT  5.110 2.740 5.360 3.480 ;
        RECT  6.720 2.620 7.000 3.480 ;
        RECT  7.760 2.620 8.040 3.480 ;
        RECT  8.800 2.620 9.080 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.260 2.600 4.250 2.760 ;
        RECT  4.090 2.160 4.250 2.760 ;
        RECT  3.260 0.460 3.420 2.760 ;
        RECT  6.960 2.300 9.440 2.460 ;
        RECT  9.280 0.860 9.440 2.460 ;
        RECT  2.840 2.300 3.420 2.460 ;
        RECT  5.840 2.280 7.120 2.440 ;
        RECT  4.090 2.160 4.630 2.320 ;
        RECT  5.840 2.000 6.000 2.440 ;
        RECT  4.470 2.000 6.000 2.160 ;
        RECT  3.140 0.460 3.420 0.680 ;
        RECT  6.260 1.810 6.480 2.120 ;
        RECT  6.260 1.810 6.740 1.970 ;
        RECT  6.580 0.810 6.740 1.970 ;
        RECT  6.580 1.340 7.140 1.620 ;
        RECT  6.320 0.810 6.740 0.970 ;
        RECT  6.320 0.440 6.480 0.970 ;
        RECT  6.200 0.440 6.480 0.660 ;
        RECT  3.580 2.180 3.930 2.440 ;
        RECT  3.580 0.460 3.740 2.440 ;
        RECT  6.080 1.260 6.360 1.580 ;
        RECT  4.220 1.260 6.360 1.420 ;
        RECT  4.220 0.460 4.380 1.420 ;
        RECT  3.580 0.460 4.380 0.620 ;
        RECT  4.980 0.940 6.060 1.100 ;
        RECT  4.980 0.460 5.140 1.100 ;
        RECT  4.540 0.460 5.140 0.740 ;
        RECT  5.520 2.600 6.060 2.760 ;
        RECT  4.500 2.480 4.950 2.640 ;
        RECT  5.520 2.340 5.680 2.760 ;
        RECT  4.790 2.340 5.680 2.500 ;
        RECT  3.900 1.580 4.300 1.980 ;
        RECT  3.900 1.580 5.880 1.740 ;
        RECT  3.900 0.840 4.060 1.980 ;
        RECT  0.600 0.560 0.760 2.190 ;
        RECT  2.940 0.880 3.100 2.080 ;
        RECT  2.820 0.560 2.980 1.040 ;
        RECT  0.600 0.560 2.980 0.720 ;
        RECT  2.460 0.880 2.620 2.320 ;
        RECT  2.460 1.380 2.780 1.660 ;
        RECT  2.400 0.880 2.620 1.160 ;
        RECT  1.240 2.150 2.240 2.310 ;
        RECT  2.080 0.920 2.240 2.310 ;
        RECT  2.080 1.460 2.300 1.740 ;
        RECT  1.240 0.920 2.240 1.080 ;
    END
END QDFFKHD

MACRO QDFFRBCHD
    CLASS CORE ;
    FOREIGN QDFFRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        RECT  6.380 1.400 6.700 1.680 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.260 1.500 1.880 ;
        RECT  1.210 1.440 1.500 1.720 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.660 8.700 2.280 ;
        RECT  8.480 2.000 8.700 2.280 ;
        RECT  8.480 0.660 8.700 0.940 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.350 -0.280 1.630 0.400 ;
        RECT  6.330 -0.280 6.610 0.400 ;
        RECT  7.900 -0.280 8.180 0.700 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.390 2.800 1.670 3.480 ;
        RECT  7.120 2.800 7.400 3.480 ;
        RECT  7.860 2.620 8.140 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.810 2.600 6.300 2.760 ;
        RECT  6.140 2.480 7.700 2.640 ;
        RECT  2.810 0.460 2.970 2.760 ;
        RECT  7.540 1.900 7.700 2.640 ;
        RECT  2.390 2.300 2.970 2.460 ;
        RECT  7.700 0.950 7.860 2.280 ;
        RECT  7.500 0.950 7.860 1.110 ;
        RECT  7.500 0.480 7.660 1.110 ;
        RECT  7.380 0.480 7.660 0.760 ;
        RECT  2.650 0.460 2.970 0.680 ;
        RECT  6.510 2.160 7.340 2.320 ;
        RECT  7.180 0.970 7.340 2.320 ;
        RECT  7.180 1.400 7.530 1.680 ;
        RECT  3.130 2.220 3.460 2.440 ;
        RECT  3.130 0.440 3.290 2.440 ;
        RECT  6.860 0.620 7.020 1.730 ;
        RECT  6.010 0.620 7.020 0.780 ;
        RECT  6.010 0.440 6.170 0.780 ;
        RECT  3.130 0.440 6.170 0.600 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.460 5.980 2.440 ;
        RECT  5.390 1.460 5.980 1.620 ;
        RECT  5.690 0.760 5.850 1.620 ;
        RECT  4.350 0.760 5.850 0.920 ;
        RECT  4.650 1.960 5.660 2.120 ;
        RECT  5.380 1.900 5.660 2.120 ;
        RECT  4.030 1.820 4.810 1.980 ;
        RECT  4.650 1.080 4.810 2.120 ;
        RECT  5.250 1.080 5.530 1.300 ;
        RECT  3.970 1.080 5.530 1.240 ;
        RECT  3.970 0.840 4.130 1.240 ;
        RECT  3.450 1.400 3.830 1.980 ;
        RECT  3.450 1.400 4.490 1.560 ;
        RECT  3.450 0.840 3.610 1.980 ;
        RECT  0.600 1.700 0.760 2.180 ;
        RECT  2.490 0.880 2.650 2.080 ;
        RECT  0.580 0.440 0.740 1.860 ;
        RECT  2.330 0.520 2.490 1.040 ;
        RECT  0.580 0.560 1.900 0.720 ;
        RECT  1.740 0.520 2.490 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.010 0.840 2.170 2.540 ;
        RECT  2.010 1.380 2.330 1.660 ;
        RECT  0.870 2.370 1.850 2.530 ;
        RECT  1.690 0.900 1.850 2.530 ;
        RECT  0.910 0.900 1.850 1.060 ;
    END
END QDFFRBCHD

MACRO QDFFRBEHD
    CLASS CORE ;
    FOREIGN QDFFRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        RECT  6.380 1.400 6.700 1.680 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.260 1.500 1.880 ;
        RECT  1.210 1.440 1.500 1.720 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.960 8.700 2.120 ;
        RECT  8.480 1.840 8.700 2.120 ;
        RECT  8.480 0.960 8.700 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.350 -0.280 1.630 0.400 ;
        RECT  6.330 -0.280 6.610 0.400 ;
        RECT  7.900 -0.280 8.180 0.580 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.390 2.800 1.670 3.480 ;
        RECT  7.170 2.800 7.450 3.480 ;
        RECT  7.900 2.620 8.180 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.810 2.600 6.300 2.760 ;
        RECT  6.140 2.480 7.700 2.640 ;
        RECT  2.810 0.460 2.970 2.760 ;
        RECT  7.540 1.900 7.700 2.640 ;
        RECT  2.390 2.300 2.970 2.460 ;
        RECT  7.700 0.960 7.860 2.280 ;
        RECT  7.540 0.960 7.860 1.240 ;
        RECT  2.650 0.460 2.970 0.680 ;
        RECT  6.560 2.160 7.340 2.320 ;
        RECT  7.180 0.480 7.340 2.320 ;
        RECT  7.180 1.400 7.540 1.680 ;
        RECT  7.180 0.480 7.400 0.760 ;
        RECT  3.130 2.220 3.460 2.440 ;
        RECT  3.130 0.440 3.290 2.440 ;
        RECT  6.860 0.620 7.020 1.730 ;
        RECT  6.010 0.620 7.020 0.780 ;
        RECT  6.010 0.440 6.170 0.780 ;
        RECT  3.130 0.440 6.170 0.600 ;
        RECT  4.400 2.280 5.980 2.440 ;
        RECT  5.820 1.460 5.980 2.440 ;
        RECT  5.390 1.460 5.980 1.620 ;
        RECT  5.690 0.760 5.850 1.620 ;
        RECT  4.350 0.760 5.850 0.920 ;
        RECT  4.650 1.960 5.660 2.120 ;
        RECT  5.380 1.900 5.660 2.120 ;
        RECT  4.030 1.820 4.810 1.980 ;
        RECT  4.650 1.080 4.810 2.120 ;
        RECT  5.250 1.080 5.530 1.300 ;
        RECT  3.970 1.080 5.530 1.240 ;
        RECT  3.970 0.840 4.130 1.240 ;
        RECT  3.450 1.400 3.830 1.980 ;
        RECT  3.450 1.400 4.490 1.560 ;
        RECT  3.450 0.840 3.610 1.980 ;
        RECT  0.600 1.700 0.760 2.180 ;
        RECT  2.490 0.880 2.650 2.080 ;
        RECT  0.580 0.440 0.740 1.860 ;
        RECT  2.330 0.520 2.490 1.040 ;
        RECT  0.580 0.560 1.900 0.720 ;
        RECT  1.740 0.520 2.490 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.010 0.840 2.170 2.540 ;
        RECT  2.010 1.380 2.330 1.660 ;
        RECT  0.870 2.360 1.850 2.520 ;
        RECT  1.690 0.900 1.850 2.520 ;
        RECT  0.910 0.900 1.850 1.060 ;
    END
END QDFFRBEHD

MACRO QDFFRBHHD
    CLASS CORE ;
    FOREIGN QDFFRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.260 1.500 1.880 ;
        RECT  1.190 1.440 1.500 1.720 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.960 9.100 2.120 ;
        RECT  8.760 1.840 9.100 2.120 ;
        RECT  8.760 0.960 9.100 1.240 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.340 -0.280 1.620 0.400 ;
        RECT  6.390 -0.280 6.670 0.400 ;
        RECT  8.180 -0.280 8.460 0.580 ;
        RECT  9.220 -0.280 9.500 0.580 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.370 2.800 1.650 3.480 ;
        RECT  6.440 2.560 6.660 3.480 ;
        RECT  7.460 2.800 7.740 3.480 ;
        RECT  8.140 2.800 8.420 3.480 ;
        RECT  9.220 2.620 9.500 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.800 2.600 6.280 2.760 ;
        RECT  6.120 2.240 6.280 2.760 ;
        RECT  2.800 0.460 2.960 2.760 ;
        RECT  2.370 2.300 2.960 2.460 ;
        RECT  6.120 2.240 8.140 2.400 ;
        RECT  7.980 0.960 8.140 2.400 ;
        RECT  7.820 1.840 8.140 2.400 ;
        RECT  7.820 0.960 8.140 1.240 ;
        RECT  2.640 0.460 2.960 0.680 ;
        RECT  6.860 1.920 7.630 2.080 ;
        RECT  7.470 0.690 7.630 2.080 ;
        RECT  7.470 1.400 7.790 1.680 ;
        RECT  7.330 0.690 7.630 0.970 ;
        RECT  3.120 2.220 3.440 2.440 ;
        RECT  3.120 0.440 3.280 2.440 ;
        RECT  6.990 1.400 7.310 1.680 ;
        RECT  6.990 0.560 7.150 1.680 ;
        RECT  6.000 0.560 7.150 0.720 ;
        RECT  3.120 0.440 6.160 0.600 ;
        RECT  4.380 2.280 5.960 2.440 ;
        RECT  5.800 1.460 5.960 2.440 ;
        RECT  5.420 1.460 5.960 1.620 ;
        RECT  5.680 0.760 5.840 1.620 ;
        RECT  4.340 0.760 5.840 0.920 ;
        RECT  4.700 1.960 5.640 2.120 ;
        RECT  5.360 1.900 5.640 2.120 ;
        RECT  4.010 1.820 4.860 1.980 ;
        RECT  4.700 1.080 4.860 2.120 ;
        RECT  5.240 1.080 5.520 1.300 ;
        RECT  3.960 1.080 5.520 1.240 ;
        RECT  3.960 0.840 4.120 1.240 ;
        RECT  3.440 1.400 3.810 1.980 ;
        RECT  3.440 1.400 4.480 1.560 ;
        RECT  3.440 0.840 3.600 1.980 ;
        RECT  0.600 1.740 0.760 2.160 ;
        RECT  2.470 0.880 2.630 2.080 ;
        RECT  0.580 0.440 0.740 1.900 ;
        RECT  2.420 0.880 2.640 1.160 ;
        RECT  2.320 0.520 2.480 1.040 ;
        RECT  0.580 0.560 1.890 0.720 ;
        RECT  1.730 0.520 2.480 0.680 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  1.990 1.950 2.150 2.540 ;
        RECT  2.000 0.840 2.160 2.110 ;
        RECT  2.000 1.380 2.310 1.660 ;
        RECT  0.860 2.370 1.830 2.530 ;
        RECT  1.670 0.910 1.830 2.530 ;
        RECT  0.900 0.910 1.830 1.070 ;
    END
END QDFFRBHHD

MACRO QDFFRBKHD
    CLASS CORE ;
    FOREIGN QDFFRBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.500 1.280 6.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.250 1.500 1.790 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.660 0.860 10.350 1.140 ;
        RECT  8.660 2.060 10.350 2.340 ;
        RECT  9.300 0.860 9.500 2.340 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 -0.280 1.780 0.400 ;
        RECT  6.510 -0.280 6.790 0.400 ;
        RECT  8.320 -0.280 8.600 0.580 ;
        RECT  9.380 -0.280 9.660 0.580 ;
        RECT  10.420 -0.280 10.700 0.580 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.500 2.800 1.780 3.480 ;
        RECT  6.570 2.560 6.790 3.480 ;
        RECT  7.590 2.800 7.870 3.480 ;
        RECT  8.340 2.560 8.620 3.480 ;
        RECT  9.380 2.620 9.660 3.480 ;
        RECT  10.420 2.620 10.700 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.920 2.600 6.410 2.760 ;
        RECT  6.250 2.240 6.410 2.760 ;
        RECT  2.920 0.460 3.080 2.760 ;
        RECT  2.500 2.300 3.080 2.460 ;
        RECT  6.250 2.240 8.300 2.400 ;
        RECT  8.140 0.890 8.300 2.400 ;
        RECT  7.980 1.840 8.300 2.400 ;
        RECT  7.980 0.960 8.300 1.240 ;
        RECT  2.760 0.460 3.080 0.680 ;
        RECT  6.990 1.920 7.750 2.080 ;
        RECT  7.590 0.960 7.750 2.080 ;
        RECT  7.590 1.400 7.950 1.680 ;
        RECT  7.450 0.960 7.750 1.240 ;
        RECT  3.240 2.220 3.570 2.440 ;
        RECT  3.240 0.440 3.400 2.440 ;
        RECT  7.110 1.400 7.430 1.680 ;
        RECT  7.110 0.560 7.270 1.680 ;
        RECT  6.120 0.560 7.270 0.720 ;
        RECT  3.240 0.440 6.280 0.600 ;
        RECT  4.510 2.280 6.090 2.440 ;
        RECT  5.930 1.460 6.090 2.440 ;
        RECT  5.530 1.460 6.090 1.620 ;
        RECT  5.800 0.760 5.960 1.620 ;
        RECT  4.460 0.760 5.960 0.920 ;
        RECT  4.820 1.960 5.770 2.120 ;
        RECT  5.490 1.900 5.770 2.120 ;
        RECT  4.140 1.820 4.980 1.980 ;
        RECT  4.820 1.080 4.980 2.120 ;
        RECT  5.360 1.080 5.640 1.300 ;
        RECT  4.080 1.080 5.640 1.240 ;
        RECT  4.080 0.840 4.240 1.240 ;
        RECT  3.560 1.400 3.940 1.980 ;
        RECT  3.560 1.400 4.640 1.560 ;
        RECT  3.560 0.840 3.720 1.980 ;
        RECT  0.600 1.720 0.760 2.180 ;
        RECT  2.600 0.880 2.760 2.080 ;
        RECT  0.580 0.440 0.740 1.880 ;
        RECT  2.440 0.560 2.600 1.040 ;
        RECT  0.580 0.560 2.600 0.720 ;
        RECT  0.580 0.440 0.860 0.720 ;
        RECT  2.120 0.880 2.280 2.540 ;
        RECT  2.120 1.380 2.440 1.660 ;
        RECT  2.060 0.880 2.280 1.160 ;
        RECT  0.900 2.420 1.900 2.580 ;
        RECT  1.740 0.910 1.900 2.580 ;
        RECT  1.740 1.440 1.960 1.720 ;
        RECT  0.900 0.910 1.900 1.070 ;
    END
END QDFFRBKHD

MACRO QDFFRSBEHD
    CLASS CORE ;
    FOREIGN QDFFRSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.770 0.840 7.100 1.340 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.420 1.500 1.700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.320 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.080 1.840 10.300 2.120 ;
        RECT  10.100 0.960 10.300 2.160 ;
        RECT  10.080 0.960 10.300 1.240 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.420 8.300 1.960 ;
        RECT  8.070 1.420 8.300 1.700 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.310 -0.280 1.590 0.400 ;
        RECT  5.430 -0.280 5.710 0.620 ;
        RECT  6.870 -0.280 7.150 0.620 ;
        RECT  8.090 -0.280 8.370 0.620 ;
        RECT  9.500 -0.280 9.780 0.580 ;
        RECT  0.000 -0.280 10.400 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.470 2.800 1.750 3.480 ;
        RECT  4.930 2.800 5.210 3.480 ;
        RECT  6.290 2.800 6.570 3.480 ;
        RECT  7.690 2.800 7.970 3.480 ;
        RECT  8.710 2.800 8.990 3.480 ;
        RECT  9.500 2.620 9.780 3.480 ;
        RECT  0.000 2.920 10.400 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.890 2.600 4.120 2.760 ;
        RECT  3.960 2.160 4.120 2.760 ;
        RECT  2.890 0.460 3.050 2.760 ;
        RECT  2.510 2.300 3.050 2.460 ;
        RECT  3.960 2.160 9.130 2.320 ;
        RECT  8.970 0.460 9.130 2.320 ;
        RECT  8.930 0.460 9.210 0.680 ;
        RECT  2.730 0.460 3.050 0.680 ;
        RECT  8.650 0.940 8.810 1.500 ;
        RECT  7.750 0.940 8.810 1.100 ;
        RECT  8.220 2.480 8.550 2.740 ;
        RECT  6.810 2.480 8.550 2.640 ;
        RECT  3.520 2.280 3.800 2.440 ;
        RECT  3.560 1.840 3.720 2.440 ;
        RECT  3.560 1.840 4.450 2.000 ;
        RECT  4.290 1.060 4.450 2.000 ;
        RECT  7.320 1.500 7.480 1.920 ;
        RECT  4.290 1.500 7.480 1.660 ;
        RECT  3.870 1.060 4.450 1.220 ;
        RECT  3.870 0.600 4.030 1.220 ;
        RECT  3.250 0.600 4.030 0.760 ;
        RECT  3.250 0.460 3.590 0.760 ;
        RECT  4.610 1.820 7.090 1.980 ;
        RECT  4.280 2.480 6.230 2.640 ;
        RECT  4.720 1.180 6.210 1.340 ;
        RECT  6.050 0.700 6.210 1.340 ;
        RECT  4.720 0.880 4.880 1.340 ;
        RECT  4.610 0.880 4.880 1.160 ;
        RECT  5.040 0.840 5.890 1.000 ;
        RECT  5.040 0.460 5.200 1.000 ;
        RECT  4.220 0.460 5.200 0.620 ;
        RECT  3.210 0.940 3.370 2.080 ;
        RECT  3.210 1.380 4.130 1.660 ;
        RECT  3.210 0.940 3.570 1.100 ;
        RECT  0.610 0.560 0.770 2.230 ;
        RECT  2.570 0.880 2.730 2.040 ;
        RECT  2.410 0.440 2.570 1.040 ;
        RECT  0.610 0.560 1.910 0.720 ;
        RECT  1.750 0.440 2.570 0.600 ;
        RECT  2.090 0.760 2.250 2.340 ;
        RECT  2.090 1.380 2.390 1.660 ;
        RECT  1.030 2.180 1.910 2.340 ;
        RECT  1.750 0.880 1.910 2.340 ;
        RECT  1.030 0.880 1.910 1.040 ;
    END
END QDFFRSBEHD

MACRO QDFFRSBHHD
    CLASS CORE ;
    FOREIGN QDFFRSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.300 1.300 7.500 2.140 ;
        RECT  7.260 1.780 7.500 2.060 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.420 1.500 1.700 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.320 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.960 0.910 10.300 2.170 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.980 8.700 1.640 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.310 -0.280 1.590 0.400 ;
        RECT  5.460 -0.280 5.680 0.680 ;
        RECT  6.980 -0.280 7.260 0.620 ;
        RECT  8.200 -0.280 8.480 0.620 ;
        RECT  9.480 -0.280 9.700 1.160 ;
        RECT  9.440 0.880 9.700 1.160 ;
        RECT  10.420 -0.280 10.700 0.580 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.470 2.800 1.750 3.480 ;
        RECT  4.930 2.800 5.210 3.480 ;
        RECT  6.350 2.800 6.630 3.480 ;
        RECT  7.110 2.800 7.390 3.480 ;
        RECT  8.310 2.800 8.590 3.480 ;
        RECT  9.340 2.800 9.620 3.480 ;
        RECT  10.420 2.620 10.700 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.890 2.600 4.120 2.760 ;
        RECT  3.960 2.160 4.120 2.760 ;
        RECT  6.420 2.480 9.800 2.640 ;
        RECT  9.640 1.320 9.800 2.640 ;
        RECT  2.890 0.460 3.050 2.760 ;
        RECT  8.870 2.240 9.150 2.640 ;
        RECT  6.420 2.160 6.580 2.640 ;
        RECT  2.510 2.300 3.050 2.460 ;
        RECT  3.960 2.160 6.580 2.320 ;
        RECT  9.120 1.320 9.800 1.480 ;
        RECT  9.120 0.460 9.280 1.480 ;
        RECT  9.000 0.460 9.320 0.720 ;
        RECT  2.730 0.460 3.050 0.680 ;
        RECT  7.670 2.160 8.340 2.320 ;
        RECT  8.180 1.000 8.340 2.320 ;
        RECT  8.180 1.850 9.370 2.010 ;
        RECT  7.980 1.000 8.340 1.160 ;
        RECT  7.980 0.840 8.140 1.160 ;
        RECT  3.520 2.280 3.800 2.440 ;
        RECT  3.560 1.840 3.720 2.440 ;
        RECT  3.560 1.840 4.450 2.000 ;
        RECT  4.290 1.060 4.450 2.000 ;
        RECT  7.860 1.320 8.020 1.940 ;
        RECT  4.290 1.500 6.770 1.660 ;
        RECT  6.610 0.900 6.770 1.660 ;
        RECT  7.660 1.320 8.020 1.480 ;
        RECT  7.660 0.900 7.820 1.480 ;
        RECT  3.870 1.060 4.450 1.220 ;
        RECT  6.610 0.900 7.820 1.060 ;
        RECT  3.870 0.600 4.030 1.220 ;
        RECT  3.250 0.600 4.030 0.760 ;
        RECT  3.250 0.460 3.590 0.760 ;
        RECT  6.750 2.100 7.090 2.320 ;
        RECT  6.750 1.820 6.910 2.320 ;
        RECT  4.610 1.820 6.910 1.980 ;
        RECT  5.040 0.840 6.000 1.000 ;
        RECT  5.840 0.560 6.000 1.000 ;
        RECT  5.040 0.460 5.200 1.000 ;
        RECT  5.840 0.560 6.600 0.720 ;
        RECT  4.220 0.460 5.200 0.620 ;
        RECT  4.720 1.180 6.380 1.340 ;
        RECT  6.160 0.880 6.380 1.340 ;
        RECT  4.720 0.880 4.880 1.340 ;
        RECT  4.610 0.880 4.880 1.160 ;
        RECT  5.530 2.480 6.190 2.760 ;
        RECT  4.280 2.480 6.190 2.640 ;
        RECT  3.210 0.940 3.370 2.080 ;
        RECT  3.210 1.380 4.130 1.660 ;
        RECT  3.210 0.940 3.570 1.100 ;
        RECT  0.610 0.560 0.770 2.230 ;
        RECT  2.570 0.880 2.730 2.040 ;
        RECT  2.410 0.440 2.570 1.040 ;
        RECT  0.610 0.560 1.910 0.720 ;
        RECT  1.750 0.440 2.570 0.600 ;
        RECT  2.090 0.760 2.250 2.340 ;
        RECT  2.090 1.380 2.390 1.660 ;
        RECT  1.030 2.180 1.910 2.340 ;
        RECT  1.750 0.880 1.910 2.340 ;
        RECT  1.030 0.880 1.910 1.040 ;
    END
END QDFFRSBHHD

MACRO QDFFSBEHD
    CLASS CORE ;
    FOREIGN QDFFSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.480 1.500 1.760 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 0.920 8.700 2.280 ;
        RECT  8.480 2.000 8.700 2.280 ;
        RECT  8.480 0.920 8.700 1.200 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.140 6.300 1.660 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.580 0.400 ;
        RECT  4.980 -0.280 5.260 0.400 ;
        RECT  7.860 -0.280 8.140 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 2.800 1.740 3.480 ;
        RECT  4.970 2.800 5.250 3.480 ;
        RECT  5.730 2.800 6.010 3.480 ;
        RECT  6.860 2.800 7.140 3.480 ;
        RECT  7.860 2.800 8.140 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.470 0.920 7.630 2.160 ;
        RECT  8.130 0.920 8.290 1.740 ;
        RECT  7.330 1.460 7.630 1.740 ;
        RECT  7.470 0.920 8.290 1.080 ;
        RECT  3.200 2.280 3.550 2.440 ;
        RECT  3.200 0.460 3.360 2.440 ;
        RECT  3.840 0.980 5.080 1.140 ;
        RECT  4.920 0.560 5.080 1.140 ;
        RECT  3.840 0.460 4.000 1.140 ;
        RECT  4.920 0.560 5.840 0.720 ;
        RECT  3.200 0.460 4.000 0.620 ;
        RECT  5.680 0.440 7.690 0.600 ;
        RECT  2.880 2.600 3.870 2.760 ;
        RECT  3.710 2.160 3.870 2.760 ;
        RECT  4.970 2.480 7.150 2.640 ;
        RECT  6.990 0.760 7.150 2.640 ;
        RECT  2.880 0.460 3.040 2.760 ;
        RECT  4.970 2.160 5.130 2.640 ;
        RECT  2.500 2.300 3.040 2.460 ;
        RECT  3.710 2.160 5.130 2.320 ;
        RECT  2.720 0.460 3.040 0.680 ;
        RECT  5.290 2.020 5.760 2.180 ;
        RECT  5.600 0.940 5.760 2.180 ;
        RECT  5.600 1.820 6.620 1.980 ;
        RECT  4.490 1.320 5.760 1.480 ;
        RECT  5.250 0.940 5.760 1.100 ;
        RECT  3.520 1.640 3.950 1.980 ;
        RECT  3.520 1.640 5.440 1.800 ;
        RECT  3.520 0.840 3.680 1.980 ;
        RECT  4.160 0.460 4.760 0.740 ;
        RECT  4.030 2.480 4.570 2.760 ;
        RECT  0.600 0.560 0.760 2.230 ;
        RECT  2.560 0.880 2.720 2.040 ;
        RECT  2.400 0.440 2.560 1.040 ;
        RECT  0.600 0.560 1.900 0.720 ;
        RECT  1.740 0.440 2.560 0.600 ;
        RECT  2.080 0.760 2.240 2.400 ;
        RECT  2.080 1.380 2.380 1.660 ;
        RECT  1.020 2.180 1.900 2.340 ;
        RECT  1.740 0.910 1.900 2.340 ;
        RECT  1.020 0.910 1.900 1.070 ;
    END
END QDFFSBEHD

MACRO QDFFSBHHD
    CLASS CORE ;
    FOREIGN QDFFSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.420 1.500 1.960 ;
        RECT  1.260 1.480 1.500 1.760 ;
        END
    END CK
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.260 0.420 1.540 ;
        RECT  0.100 1.090 0.300 1.630 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.740 9.100 2.460 ;
        RECT  8.700 2.300 9.100 2.460 ;
        RECT  8.760 0.740 9.100 1.020 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 1.140 6.300 1.660 ;
        END
    END SB
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.300 -0.280 1.580 0.400 ;
        RECT  4.920 -0.280 5.200 0.400 ;
        RECT  6.190 -0.280 6.470 0.400 ;
        RECT  8.140 -0.280 8.420 0.400 ;
        RECT  9.220 -0.280 9.500 0.580 ;
        RECT  0.000 -0.280 9.600 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.460 2.800 1.740 3.480 ;
        RECT  5.010 2.800 5.290 3.480 ;
        RECT  6.150 2.800 6.430 3.480 ;
        RECT  7.270 2.800 7.550 3.480 ;
        RECT  8.180 2.620 8.460 3.480 ;
        RECT  9.220 2.620 9.500 3.480 ;
        RECT  0.000 2.920 9.600 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  7.610 1.900 8.680 2.060 ;
        RECT  8.520 1.400 8.680 2.060 ;
        RECT  7.610 0.960 7.770 2.060 ;
        RECT  7.500 1.340 7.770 1.620 ;
        RECT  3.200 2.280 3.550 2.440 ;
        RECT  3.200 0.460 3.360 2.440 ;
        RECT  8.040 0.560 8.200 1.620 ;
        RECT  3.840 0.880 5.210 1.040 ;
        RECT  5.050 0.560 5.210 1.040 ;
        RECT  3.840 0.460 4.000 1.040 ;
        RECT  5.050 0.560 8.200 0.720 ;
        RECT  3.200 0.460 4.000 0.620 ;
        RECT  2.880 2.600 3.870 2.760 ;
        RECT  3.710 2.160 3.870 2.760 ;
        RECT  4.990 2.480 7.080 2.640 ;
        RECT  6.920 1.020 7.080 2.640 ;
        RECT  2.880 0.460 3.040 2.760 ;
        RECT  6.770 2.320 7.080 2.640 ;
        RECT  4.990 2.160 5.150 2.640 ;
        RECT  2.500 2.300 3.040 2.460 ;
        RECT  3.710 2.160 5.150 2.320 ;
        RECT  6.920 1.020 7.350 1.180 ;
        RECT  2.720 0.460 3.040 0.680 ;
        RECT  5.570 0.880 5.730 2.210 ;
        RECT  4.470 1.200 4.750 1.660 ;
        RECT  4.470 1.200 5.730 1.360 ;
        RECT  5.370 0.880 5.730 1.360 ;
        RECT  3.520 1.820 5.390 1.980 ;
        RECT  5.110 1.520 5.390 1.980 ;
        RECT  3.520 0.840 3.680 1.980 ;
        RECT  4.250 2.480 4.790 2.760 ;
        RECT  4.160 0.440 4.760 0.720 ;
        RECT  0.600 0.560 0.760 2.230 ;
        RECT  2.560 0.880 2.720 2.040 ;
        RECT  2.400 0.440 2.560 1.040 ;
        RECT  0.600 0.560 1.900 0.720 ;
        RECT  1.740 0.440 2.560 0.600 ;
        RECT  2.080 0.760 2.240 2.400 ;
        RECT  2.080 1.380 2.380 1.660 ;
        RECT  1.020 2.180 1.900 2.340 ;
        RECT  1.740 0.910 1.900 2.340 ;
        RECT  1.020 0.910 1.900 1.070 ;
    END
END QDFFSBHHD

MACRO QDFZCHD
    CLASS CORE ;
    FOREIGN QDFZCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.310 3.190 1.590 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 0.440 9.900 2.120 ;
        RECT  9.680 1.840 9.900 2.120 ;
        RECT  9.620 0.440 9.900 0.660 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 3.420 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  8.180 -0.280 8.460 0.420 ;
        RECT  9.000 -0.280 9.280 0.600 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.520 3.480 ;
        RECT  6.570 2.800 6.850 3.480 ;
        RECT  7.620 2.800 8.360 3.480 ;
        RECT  9.000 2.060 9.280 2.280 ;
        RECT  9.080 2.060 9.280 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.580 2.540 8.920 2.760 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  7.710 2.480 8.740 2.640 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  8.580 0.860 8.740 2.760 ;
        RECT  7.710 1.860 7.870 2.640 ;
        RECT  4.240 2.300 4.820 2.460 ;
        RECT  5.490 2.160 6.030 2.320 ;
        RECT  5.870 1.860 6.030 2.320 ;
        RECT  5.870 1.860 7.870 2.020 ;
        RECT  8.570 0.860 8.900 1.080 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  8.120 0.580 8.280 2.120 ;
        RECT  8.120 1.340 8.420 1.620 ;
        RECT  7.580 0.580 8.280 0.740 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.780 1.140 7.940 1.660 ;
        RECT  5.620 1.140 7.940 1.300 ;
        RECT  5.620 0.460 5.780 1.300 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  7.140 0.580 7.420 0.980 ;
        RECT  5.940 0.580 7.420 0.740 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  5.900 2.480 6.430 2.640 ;
        RECT  7.140 2.180 7.420 2.520 ;
        RECT  6.270 2.360 7.420 2.520 ;
        RECT  5.300 1.460 5.700 1.980 ;
        RECT  5.300 1.460 7.280 1.620 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.660 0.560 3.740 0.720 ;
        RECT  3.580 0.440 4.380 0.600 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  3.860 0.840 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.920 3.680 2.310 ;
        RECT  2.760 0.920 3.680 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END QDFZCHD

MACRO QDFZEHD
    CLASS CORE ;
    FOREIGN QDFZEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.350 3.190 1.630 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.300 0.440 9.500 2.120 ;
        RECT  9.140 1.840 9.500 2.120 ;
        RECT  9.080 0.440 9.500 0.660 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 3.330 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  8.180 -0.280 8.460 0.420 ;
        RECT  9.660 -0.280 9.880 0.660 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.520 3.480 ;
        RECT  6.570 2.800 6.850 3.480 ;
        RECT  7.620 2.800 8.360 3.480 ;
        RECT  9.600 2.620 9.880 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  8.580 2.540 8.920 2.760 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  7.710 2.480 8.740 2.640 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  8.580 0.860 8.740 2.760 ;
        RECT  7.710 1.860 7.870 2.640 ;
        RECT  4.240 2.300 4.820 2.460 ;
        RECT  5.490 2.160 6.030 2.320 ;
        RECT  5.870 1.860 6.030 2.320 ;
        RECT  5.870 1.860 7.870 2.020 ;
        RECT  8.570 0.860 8.900 1.080 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  8.120 0.580 8.280 2.080 ;
        RECT  8.120 1.340 8.420 1.620 ;
        RECT  7.580 0.580 8.280 0.740 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.780 1.140 7.940 1.660 ;
        RECT  5.620 1.140 7.940 1.300 ;
        RECT  5.620 0.460 5.780 1.300 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  7.140 0.580 7.420 0.980 ;
        RECT  5.940 0.580 7.420 0.740 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  5.900 2.480 6.430 2.640 ;
        RECT  7.140 2.180 7.420 2.520 ;
        RECT  6.270 2.360 7.420 2.520 ;
        RECT  5.300 1.460 5.700 1.980 ;
        RECT  5.300 1.460 7.280 1.620 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.660 0.560 3.680 0.720 ;
        RECT  3.520 0.440 4.380 0.600 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  3.860 0.760 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.920 3.680 2.310 ;
        RECT  2.760 0.920 3.680 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END QDFZEHD

MACRO QDFZHHD
    CLASS CORE ;
    FOREIGN QDFZHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.350 3.190 1.630 ;
        RECT  2.900 1.240 3.100 1.780 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.880 9.100 2.120 ;
        RECT  8.640 1.840 9.100 2.120 ;
        RECT  8.640 0.880 9.100 1.160 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 3.330 0.400 ;
        RECT  6.700 -0.280 6.980 0.420 ;
        RECT  8.060 -0.280 8.340 0.580 ;
        RECT  9.100 -0.280 9.380 0.580 ;
        RECT  0.000 -0.280 10.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.520 3.480 ;
        RECT  6.490 2.800 6.770 3.480 ;
        RECT  8.060 2.620 8.340 3.480 ;
        RECT  9.100 2.620 9.380 3.480 ;
        RECT  0.000 2.920 10.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.660 2.600 5.650 2.760 ;
        RECT  5.490 2.160 5.650 2.760 ;
        RECT  4.660 0.460 4.820 2.760 ;
        RECT  7.620 2.300 9.840 2.460 ;
        RECT  9.680 0.910 9.840 2.460 ;
        RECT  4.240 2.300 4.820 2.460 ;
        RECT  7.220 2.220 7.780 2.380 ;
        RECT  5.490 2.160 6.030 2.320 ;
        RECT  7.220 2.030 7.380 2.380 ;
        RECT  5.870 2.030 7.380 2.190 ;
        RECT  4.540 0.460 4.820 0.680 ;
        RECT  7.540 1.840 8.070 2.060 ;
        RECT  7.910 1.000 8.070 2.060 ;
        RECT  7.910 1.340 8.480 1.620 ;
        RECT  7.700 1.000 8.070 1.160 ;
        RECT  7.700 0.440 7.860 1.160 ;
        RECT  7.500 0.440 7.860 0.600 ;
        RECT  4.980 2.180 5.330 2.440 ;
        RECT  4.980 0.460 5.140 2.440 ;
        RECT  7.490 1.350 7.710 1.630 ;
        RECT  5.620 1.350 7.710 1.510 ;
        RECT  5.620 0.460 5.780 1.510 ;
        RECT  4.980 0.460 5.780 0.620 ;
        RECT  6.380 0.940 7.460 1.100 ;
        RECT  6.380 0.460 6.540 1.100 ;
        RECT  5.940 0.460 6.540 0.740 ;
        RECT  6.900 2.540 7.460 2.700 ;
        RECT  5.900 2.480 6.430 2.640 ;
        RECT  6.900 2.360 7.060 2.700 ;
        RECT  6.270 2.360 7.060 2.520 ;
        RECT  5.300 1.680 5.700 1.980 ;
        RECT  5.300 1.680 7.280 1.840 ;
        RECT  5.300 0.840 5.460 1.980 ;
        RECT  1.480 2.600 2.300 2.760 ;
        RECT  2.140 0.560 2.300 2.760 ;
        RECT  4.340 0.880 4.500 2.080 ;
        RECT  4.220 0.440 4.380 1.040 ;
        RECT  1.660 0.560 3.680 0.720 ;
        RECT  3.520 0.440 4.380 0.600 ;
        RECT  1.660 0.460 1.940 0.720 ;
        RECT  3.860 0.760 4.020 2.320 ;
        RECT  3.860 1.380 4.160 1.660 ;
        RECT  2.760 2.150 3.680 2.310 ;
        RECT  3.520 0.920 3.680 2.310 ;
        RECT  2.760 0.920 3.680 1.080 ;
        RECT  1.760 2.140 1.980 2.420 ;
        RECT  0.920 2.200 1.980 2.360 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 0.800 1.080 2.360 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END QDFZHHD

MACRO QDFZKHD
    CLASS CORE ;
    FOREIGN QDFZKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.240 3.500 1.780 ;
        RECT  3.260 1.350 3.500 1.630 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.250 2.700 1.780 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 0.880 10.100 1.160 ;
        RECT  8.900 1.840 10.100 2.120 ;
        RECT  9.300 0.880 9.500 2.120 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.440 -0.280 3.720 0.400 ;
        RECT  6.900 -0.280 7.180 0.420 ;
        RECT  8.320 -0.280 8.600 0.580 ;
        RECT  9.360 -0.280 9.640 0.580 ;
        RECT  10.400 -0.280 10.680 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 3.720 3.480 ;
        RECT  6.740 2.800 7.020 3.480 ;
        RECT  8.320 2.620 8.600 3.480 ;
        RECT  9.360 2.620 9.640 3.480 ;
        RECT  10.400 2.620 10.680 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.860 2.600 5.850 2.760 ;
        RECT  5.690 2.160 5.850 2.760 ;
        RECT  4.860 0.460 5.020 2.760 ;
        RECT  8.560 2.300 11.040 2.460 ;
        RECT  10.880 0.860 11.040 2.460 ;
        RECT  4.440 2.300 5.020 2.460 ;
        RECT  7.500 2.280 8.720 2.440 ;
        RECT  5.690 2.160 6.230 2.320 ;
        RECT  7.500 2.000 7.660 2.440 ;
        RECT  6.070 2.000 7.660 2.160 ;
        RECT  4.740 0.460 5.020 0.680 ;
        RECT  7.860 1.810 8.080 2.120 ;
        RECT  7.860 1.810 8.340 1.970 ;
        RECT  8.180 0.810 8.340 1.970 ;
        RECT  8.180 1.340 8.740 1.620 ;
        RECT  7.920 0.810 8.340 0.970 ;
        RECT  7.920 0.440 8.080 0.970 ;
        RECT  7.800 0.440 8.080 0.660 ;
        RECT  5.180 2.180 5.530 2.440 ;
        RECT  5.180 0.460 5.340 2.440 ;
        RECT  7.680 1.260 7.960 1.580 ;
        RECT  5.820 1.260 7.960 1.420 ;
        RECT  5.820 0.460 5.980 1.420 ;
        RECT  5.180 0.460 5.980 0.620 ;
        RECT  6.580 0.940 7.660 1.100 ;
        RECT  6.580 0.460 6.740 1.100 ;
        RECT  6.140 0.460 6.740 0.740 ;
        RECT  7.180 2.600 7.660 2.760 ;
        RECT  6.100 2.480 6.630 2.640 ;
        RECT  7.180 2.340 7.340 2.760 ;
        RECT  6.470 2.340 7.340 2.500 ;
        RECT  5.500 1.580 5.900 1.980 ;
        RECT  5.500 1.580 7.480 1.740 ;
        RECT  5.500 0.840 5.660 1.980 ;
        RECT  1.480 2.380 2.300 2.540 ;
        RECT  2.140 0.460 2.300 2.540 ;
        RECT  4.540 0.880 4.700 2.080 ;
        RECT  4.420 0.560 4.580 1.040 ;
        RECT  2.140 0.560 4.580 0.720 ;
        RECT  1.620 0.460 2.300 0.620 ;
        RECT  4.060 0.880 4.220 2.320 ;
        RECT  4.060 1.380 4.380 1.660 ;
        RECT  4.000 0.880 4.220 1.160 ;
        RECT  2.840 2.150 3.840 2.310 ;
        RECT  3.680 0.920 3.840 2.310 ;
        RECT  3.680 1.460 3.900 1.740 ;
        RECT  2.840 0.920 3.840 1.080 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.920 2.060 1.980 2.220 ;
        RECT  1.760 1.940 1.980 2.220 ;
        RECT  0.920 0.800 1.080 2.220 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  0.100 0.460 0.380 1.040 ;
        RECT  0.100 0.800 1.080 0.960 ;
    END
END QDFZKHD

MACRO QDFZRBCHD
    CLASS CORE ;
    FOREIGN QDFZRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.530 11.100 2.640 ;
        RECT  10.880 2.360 11.100 2.640 ;
        RECT  10.880 0.650 11.100 0.930 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.540 -0.280 3.820 0.400 ;
        RECT  8.520 -0.280 8.740 0.500 ;
        RECT  10.260 -0.280 10.540 0.400 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.560 2.800 3.840 3.480 ;
        RECT  8.040 2.800 8.720 3.480 ;
        RECT  9.560 2.800 9.840 3.480 ;
        RECT  10.260 2.800 10.540 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.000 2.600 6.080 2.760 ;
        RECT  5.920 2.140 6.080 2.760 ;
        RECT  7.800 2.480 10.180 2.640 ;
        RECT  10.020 0.800 10.180 2.640 ;
        RECT  5.000 0.460 5.160 2.760 ;
        RECT  7.800 2.140 7.960 2.640 ;
        RECT  4.580 2.300 5.160 2.460 ;
        RECT  5.920 2.140 7.960 2.300 ;
        RECT  9.780 0.800 10.180 0.960 ;
        RECT  4.840 0.460 5.160 0.680 ;
        RECT  8.960 2.160 9.860 2.320 ;
        RECT  9.700 1.120 9.860 2.320 ;
        RECT  9.380 1.120 9.860 1.280 ;
        RECT  9.380 0.920 9.540 1.280 ;
        RECT  5.320 2.220 5.650 2.440 ;
        RECT  5.320 0.440 5.480 2.440 ;
        RECT  8.920 1.460 9.490 1.620 ;
        RECT  8.920 0.660 9.080 1.620 ;
        RECT  8.200 0.660 9.080 0.820 ;
        RECT  8.200 0.440 8.360 0.820 ;
        RECT  5.320 0.440 8.360 0.600 ;
        RECT  8.120 1.820 8.280 2.220 ;
        RECT  6.220 1.820 8.280 1.980 ;
        RECT  7.270 1.080 7.430 1.980 ;
        RECT  7.270 1.080 7.720 1.300 ;
        RECT  6.160 1.080 7.720 1.240 ;
        RECT  6.160 0.840 6.320 1.240 ;
        RECT  7.600 1.460 8.040 1.620 ;
        RECT  7.880 0.760 8.040 1.620 ;
        RECT  6.540 0.760 8.040 0.920 ;
        RECT  7.420 2.460 7.640 2.740 ;
        RECT  6.500 2.460 7.640 2.620 ;
        RECT  5.640 1.400 6.020 1.980 ;
        RECT  5.640 1.400 7.100 1.560 ;
        RECT  5.640 0.840 5.800 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.680 0.880 4.840 2.080 ;
        RECT  4.520 0.520 4.680 1.040 ;
        RECT  1.620 0.560 4.090 0.720 ;
        RECT  3.930 0.520 4.680 0.680 ;
        RECT  4.200 0.840 4.360 2.540 ;
        RECT  4.200 1.380 4.520 1.660 ;
        RECT  2.940 2.320 4.040 2.480 ;
        RECT  3.880 0.880 4.040 2.480 ;
        RECT  2.940 0.880 4.040 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END QDFZRBCHD

MACRO QDFZRBEHD
    CLASS CORE ;
    FOREIGN QDFZRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.440 3.560 1.720 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.700 2.120 ;
        RECT  10.360 1.840 10.700 2.120 ;
        RECT  10.360 0.960 10.700 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.560 -0.280 3.840 0.400 ;
        RECT  8.540 -0.280 8.820 0.400 ;
        RECT  9.400 -0.280 9.680 0.400 ;
        RECT  10.820 -0.280 11.100 0.580 ;
        RECT  0.000 -0.280 11.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.580 2.800 3.860 3.480 ;
        RECT  9.430 2.800 9.710 3.480 ;
        RECT  10.820 2.620 11.100 3.480 ;
        RECT  0.000 2.920 11.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.020 2.600 8.510 2.760 ;
        RECT  10.020 0.440 10.180 2.640 ;
        RECT  8.350 2.480 10.180 2.640 ;
        RECT  5.020 0.460 5.180 2.760 ;
        RECT  4.600 2.300 5.180 2.460 ;
        RECT  9.960 0.440 10.180 0.720 ;
        RECT  4.860 0.460 5.180 0.680 ;
        RECT  8.820 2.160 9.550 2.320 ;
        RECT  9.390 0.970 9.550 2.320 ;
        RECT  9.390 1.460 9.750 1.740 ;
        RECT  5.340 2.220 5.670 2.440 ;
        RECT  5.340 0.440 5.500 2.440 ;
        RECT  9.070 0.620 9.230 1.730 ;
        RECT  8.220 0.620 9.230 0.780 ;
        RECT  8.220 0.440 8.380 0.780 ;
        RECT  5.340 0.440 8.380 0.600 ;
        RECT  6.610 2.280 8.190 2.440 ;
        RECT  8.030 1.460 8.190 2.440 ;
        RECT  7.600 1.460 8.190 1.620 ;
        RECT  7.900 0.760 8.060 1.620 ;
        RECT  6.560 0.760 8.060 0.920 ;
        RECT  6.860 1.960 7.870 2.120 ;
        RECT  7.590 1.900 7.870 2.120 ;
        RECT  6.240 1.820 7.020 1.980 ;
        RECT  6.860 1.080 7.020 2.120 ;
        RECT  7.460 1.080 7.740 1.300 ;
        RECT  6.180 1.080 7.740 1.240 ;
        RECT  6.180 0.840 6.340 1.240 ;
        RECT  5.660 1.400 6.040 1.980 ;
        RECT  5.660 1.400 6.700 1.560 ;
        RECT  5.660 0.840 5.820 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.700 0.880 4.860 2.080 ;
        RECT  4.540 0.520 4.700 1.040 ;
        RECT  1.620 0.560 4.110 0.720 ;
        RECT  3.950 0.520 4.700 0.680 ;
        RECT  4.220 0.840 4.380 2.540 ;
        RECT  4.220 1.380 4.540 1.660 ;
        RECT  2.960 2.420 4.060 2.580 ;
        RECT  3.900 0.880 4.060 2.580 ;
        RECT  2.960 0.880 4.060 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END QDFZRBEHD

MACRO QDFZRBHHD
    CLASS CORE ;
    FOREIGN QDFZRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.440 3.560 1.720 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 0.960 11.500 2.120 ;
        RECT  11.160 1.840 11.500 2.120 ;
        RECT  11.160 0.960 11.500 1.240 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.560 -0.280 3.840 0.400 ;
        RECT  8.610 -0.280 8.890 0.400 ;
        RECT  10.580 -0.280 10.860 0.580 ;
        RECT  11.620 -0.280 11.900 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.580 2.800 3.860 3.480 ;
        RECT  8.670 2.740 10.010 3.480 ;
        RECT  10.540 2.800 10.820 3.480 ;
        RECT  11.620 2.620 11.900 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.020 2.600 8.510 2.760 ;
        RECT  8.350 2.420 8.510 2.760 ;
        RECT  5.020 0.460 5.180 2.760 ;
        RECT  8.350 2.420 10.380 2.580 ;
        RECT  10.220 0.890 10.380 2.580 ;
        RECT  4.600 2.300 5.180 2.460 ;
        RECT  4.860 0.460 5.180 0.680 ;
        RECT  9.130 2.100 9.850 2.260 ;
        RECT  9.690 0.600 9.850 2.260 ;
        RECT  9.690 1.460 10.050 1.740 ;
        RECT  5.340 2.220 5.670 2.440 ;
        RECT  5.340 0.440 5.500 2.440 ;
        RECT  9.370 0.560 9.530 1.680 ;
        RECT  8.220 0.560 9.530 0.720 ;
        RECT  5.340 0.440 8.380 0.600 ;
        RECT  6.610 2.280 8.190 2.440 ;
        RECT  8.030 1.460 8.190 2.440 ;
        RECT  7.640 1.460 8.190 1.620 ;
        RECT  7.900 0.760 8.060 1.620 ;
        RECT  6.560 0.760 8.060 0.920 ;
        RECT  6.920 1.960 7.870 2.120 ;
        RECT  7.590 1.900 7.870 2.120 ;
        RECT  6.240 1.820 7.080 1.980 ;
        RECT  6.920 1.080 7.080 2.120 ;
        RECT  7.460 1.080 7.740 1.300 ;
        RECT  6.180 1.080 7.740 1.240 ;
        RECT  6.180 0.840 6.340 1.240 ;
        RECT  5.660 1.400 6.040 1.980 ;
        RECT  5.660 1.400 6.700 1.560 ;
        RECT  5.660 0.840 5.820 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.700 0.880 4.860 2.080 ;
        RECT  4.540 0.520 4.700 1.040 ;
        RECT  1.620 0.560 4.110 0.720 ;
        RECT  3.950 0.520 4.700 0.680 ;
        RECT  4.220 0.840 4.380 2.540 ;
        RECT  4.220 1.380 4.540 1.660 ;
        RECT  2.960 2.420 4.060 2.580 ;
        RECT  3.900 0.880 4.060 2.580 ;
        RECT  2.960 0.880 4.060 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END QDFZRBHHD

MACRO QDFZRBKHD
    CLASS CORE ;
    FOREIGN QDFZRBKHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.500 1.280 8.700 1.940 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.440 3.560 1.720 ;
        RECT  3.300 1.200 3.500 1.740 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.200 3.100 1.800 ;
        RECT  2.740 1.340 3.100 1.620 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.560 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.060 0.860 12.750 1.140 ;
        RECT  11.060 2.060 12.750 2.340 ;
        RECT  11.700 0.860 11.900 2.340 ;
        END
    END Q
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.540 -0.280 2.820 0.400 ;
        RECT  3.560 -0.280 3.840 0.400 ;
        RECT  8.610 -0.280 8.890 0.400 ;
        RECT  10.720 -0.280 11.000 0.580 ;
        RECT  11.780 -0.280 12.060 0.580 ;
        RECT  12.820 -0.280 13.100 0.580 ;
        RECT  0.000 -0.280 13.200 0.280 ;
        RECT  0.620 -0.280 0.900 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.580 2.800 3.860 3.480 ;
        RECT  8.670 2.740 10.010 3.480 ;
        RECT  10.700 2.800 10.980 3.480 ;
        RECT  11.780 2.620 12.060 3.480 ;
        RECT  12.820 2.620 13.100 3.480 ;
        RECT  0.000 2.920 13.200 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.020 2.600 8.510 2.760 ;
        RECT  8.350 2.420 8.510 2.760 ;
        RECT  5.020 0.460 5.180 2.760 ;
        RECT  8.350 2.420 10.380 2.580 ;
        RECT  10.220 0.890 10.380 2.580 ;
        RECT  4.600 2.300 5.180 2.460 ;
        RECT  4.860 0.460 5.180 0.680 ;
        RECT  9.130 2.100 9.850 2.260 ;
        RECT  9.690 0.600 9.850 2.260 ;
        RECT  9.690 1.460 10.050 1.740 ;
        RECT  5.340 2.220 5.670 2.440 ;
        RECT  5.340 0.440 5.500 2.440 ;
        RECT  9.370 0.560 9.530 1.680 ;
        RECT  8.220 0.560 9.530 0.720 ;
        RECT  5.340 0.440 8.380 0.600 ;
        RECT  6.610 2.280 8.190 2.440 ;
        RECT  8.030 1.460 8.190 2.440 ;
        RECT  7.630 1.460 8.190 1.620 ;
        RECT  7.900 0.760 8.060 1.620 ;
        RECT  6.560 0.760 8.060 0.920 ;
        RECT  6.920 1.960 7.870 2.120 ;
        RECT  7.590 1.900 7.870 2.120 ;
        RECT  6.240 1.820 7.080 1.980 ;
        RECT  6.920 1.080 7.080 2.120 ;
        RECT  7.460 1.080 7.740 1.300 ;
        RECT  6.180 1.080 7.740 1.240 ;
        RECT  6.180 0.840 6.340 1.240 ;
        RECT  5.660 1.400 6.040 1.980 ;
        RECT  5.660 1.400 6.740 1.560 ;
        RECT  5.660 0.840 5.820 1.980 ;
        RECT  1.520 2.520 2.360 2.680 ;
        RECT  2.200 0.560 2.360 2.680 ;
        RECT  4.700 0.880 4.860 2.080 ;
        RECT  4.540 0.520 4.700 1.040 ;
        RECT  1.620 0.560 4.110 0.720 ;
        RECT  3.950 0.520 4.700 0.680 ;
        RECT  4.220 0.840 4.380 2.540 ;
        RECT  4.220 1.380 4.540 1.660 ;
        RECT  2.960 2.420 4.060 2.580 ;
        RECT  3.900 0.880 4.060 2.580 ;
        RECT  2.960 0.880 4.060 1.040 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.460 0.260 2.280 ;
        RECT  1.880 0.880 2.040 1.780 ;
        RECT  0.920 0.880 1.080 1.460 ;
        RECT  0.100 0.880 2.040 1.040 ;
        RECT  0.100 0.460 0.380 1.040 ;
    END
END QDFZRBKHD

MACRO QDFZRSBEHD
    CLASS CORE ;
    FOREIGN QDFZRSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.780 0.840 9.100 1.340 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.110 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.420 2.300 1.990 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.960 11.260 1.240 ;
        RECT  10.900 1.840 11.260 2.120 ;
        RECT  10.900 0.960 11.100 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  9.700 1.420 9.920 1.700 ;
        RECT  9.700 1.420 9.900 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 -0.280 3.280 0.400 ;
        RECT  7.120 -0.280 7.400 0.620 ;
        RECT  8.560 -0.280 8.840 0.620 ;
        RECT  9.780 -0.280 10.060 0.620 ;
        RECT  11.500 -0.280 11.780 0.580 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 2.800 2.620 3.480 ;
        RECT  3.160 2.800 3.440 3.480 ;
        RECT  6.620 2.800 6.900 3.480 ;
        RECT  8.220 2.800 8.500 3.480 ;
        RECT  9.380 2.800 9.660 3.480 ;
        RECT  10.400 2.800 10.680 3.480 ;
        RECT  11.500 2.620 11.780 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.560 2.620 0.840 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.580 2.600 5.810 2.760 ;
        RECT  5.650 2.160 5.810 2.760 ;
        RECT  4.580 0.460 4.740 2.760 ;
        RECT  4.200 2.300 4.740 2.460 ;
        RECT  5.650 2.160 10.740 2.320 ;
        RECT  10.580 0.460 10.740 2.320 ;
        RECT  10.580 0.460 10.900 0.680 ;
        RECT  4.420 0.460 4.740 0.680 ;
        RECT  10.240 0.940 10.400 1.460 ;
        RECT  9.440 0.940 10.400 1.100 ;
        RECT  9.910 2.480 10.240 2.740 ;
        RECT  8.740 2.480 10.240 2.640 ;
        RECT  5.210 2.280 5.490 2.440 ;
        RECT  5.250 1.840 5.410 2.440 ;
        RECT  5.250 1.840 6.140 2.000 ;
        RECT  5.980 1.060 6.140 2.000 ;
        RECT  9.180 1.500 9.340 1.920 ;
        RECT  5.980 1.500 9.340 1.660 ;
        RECT  5.560 1.060 6.140 1.220 ;
        RECT  5.560 0.600 5.720 1.220 ;
        RECT  4.940 0.600 5.720 0.760 ;
        RECT  4.940 0.460 5.280 0.760 ;
        RECT  6.300 1.820 9.020 1.980 ;
        RECT  5.970 2.480 8.160 2.640 ;
        RECT  6.410 1.180 7.900 1.340 ;
        RECT  7.740 0.700 7.900 1.340 ;
        RECT  6.410 0.880 6.570 1.340 ;
        RECT  6.300 0.880 6.570 1.160 ;
        RECT  6.730 0.840 7.580 1.000 ;
        RECT  6.730 0.460 6.890 1.000 ;
        RECT  5.910 0.460 6.890 0.620 ;
        RECT  4.900 0.940 5.060 2.080 ;
        RECT  4.900 1.380 5.820 1.660 ;
        RECT  4.900 0.940 5.260 1.100 ;
        RECT  1.360 2.220 1.880 2.380 ;
        RECT  1.720 0.460 1.880 2.380 ;
        RECT  4.260 0.880 4.420 2.040 ;
        RECT  4.100 0.440 4.260 1.040 ;
        RECT  1.720 0.560 3.600 0.720 ;
        RECT  1.640 0.460 1.960 0.620 ;
        RECT  3.440 0.440 4.260 0.600 ;
        RECT  3.780 0.760 3.940 2.340 ;
        RECT  3.780 1.380 4.080 1.660 ;
        RECT  2.680 2.240 3.600 2.400 ;
        RECT  3.440 0.940 3.600 2.400 ;
        RECT  2.680 0.940 3.600 1.100 ;
        RECT  1.020 2.600 1.960 2.760 ;
        RECT  1.020 2.200 1.180 2.760 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END QDFZRSBEHD

MACRO QDFZRSBHHD
    CLASS CORE ;
    FOREIGN QDFZRSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.900 1.780 9.130 2.060 ;
        RECT  8.900 1.640 9.100 2.140 ;
        END
    END RB
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.420 3.110 1.700 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.420 2.300 1.990 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.900 0.960 12.300 2.120 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.100 1.420 10.390 1.700 ;
        RECT  10.100 1.420 10.300 1.960 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.560 -0.280 2.840 0.400 ;
        RECT  3.000 -0.280 3.280 0.400 ;
        RECT  7.170 -0.280 7.390 0.680 ;
        RECT  8.690 -0.280 8.970 0.620 ;
        RECT  10.010 -0.280 10.290 0.660 ;
        RECT  11.340 -0.280 11.620 0.400 ;
        RECT  12.420 -0.280 12.700 0.580 ;
        RECT  0.000 -0.280 12.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.340 2.800 2.620 3.480 ;
        RECT  3.160 2.800 3.440 3.480 ;
        RECT  6.620 2.800 6.900 3.480 ;
        RECT  8.040 2.800 8.320 3.480 ;
        RECT  8.870 2.800 9.150 3.480 ;
        RECT  10.070 2.800 10.350 3.480 ;
        RECT  11.340 2.800 11.620 3.480 ;
        RECT  12.420 2.620 12.700 3.480 ;
        RECT  0.000 2.920 12.800 3.480 ;
        RECT  0.560 2.620 0.840 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.580 2.600 5.810 2.760 ;
        RECT  5.650 2.160 5.810 2.760 ;
        RECT  7.980 2.480 11.500 2.640 ;
        RECT  11.340 0.590 11.500 2.640 ;
        RECT  4.580 0.460 4.740 2.760 ;
        RECT  7.980 2.160 8.140 2.640 ;
        RECT  4.200 2.300 4.740 2.460 ;
        RECT  5.650 2.160 8.140 2.320 ;
        RECT  10.910 0.590 11.500 0.750 ;
        RECT  4.420 0.460 4.740 0.680 ;
        RECT  10.910 0.440 11.130 0.750 ;
        RECT  9.430 2.160 11.170 2.320 ;
        RECT  11.010 1.240 11.170 2.320 ;
        RECT  10.570 1.240 11.170 1.400 ;
        RECT  10.570 0.870 10.730 1.400 ;
        RECT  9.630 0.780 9.850 1.140 ;
        RECT  9.630 0.870 10.730 1.030 ;
        RECT  5.210 2.280 5.490 2.440 ;
        RECT  5.250 1.840 5.410 2.440 ;
        RECT  5.250 1.840 6.140 2.000 ;
        RECT  5.980 1.060 6.140 2.000 ;
        RECT  9.750 1.300 9.910 1.940 ;
        RECT  5.980 1.500 8.460 1.660 ;
        RECT  8.300 0.900 8.460 1.660 ;
        RECT  9.310 1.300 9.910 1.460 ;
        RECT  9.310 0.900 9.470 1.460 ;
        RECT  5.560 1.060 6.140 1.220 ;
        RECT  8.300 0.900 9.470 1.060 ;
        RECT  5.560 0.600 5.720 1.220 ;
        RECT  4.940 0.600 5.720 0.760 ;
        RECT  4.940 0.460 5.280 0.760 ;
        RECT  8.400 1.820 8.740 2.320 ;
        RECT  6.300 1.820 8.740 1.980 ;
        RECT  6.730 0.840 7.710 1.000 ;
        RECT  7.550 0.560 7.710 1.000 ;
        RECT  6.730 0.460 6.890 1.000 ;
        RECT  7.550 0.560 8.270 0.720 ;
        RECT  5.910 0.460 6.890 0.620 ;
        RECT  6.410 1.180 8.090 1.340 ;
        RECT  7.870 0.880 8.090 1.340 ;
        RECT  6.410 0.880 6.570 1.340 ;
        RECT  6.300 0.880 6.570 1.160 ;
        RECT  7.220 2.480 7.820 2.760 ;
        RECT  5.970 2.480 7.820 2.640 ;
        RECT  4.900 0.940 5.060 2.080 ;
        RECT  4.900 1.380 5.820 1.660 ;
        RECT  4.900 0.940 5.260 1.100 ;
        RECT  1.360 2.220 1.880 2.380 ;
        RECT  1.720 0.460 1.880 2.380 ;
        RECT  4.260 0.880 4.420 2.040 ;
        RECT  4.100 0.440 4.260 1.040 ;
        RECT  1.720 0.560 3.600 0.720 ;
        RECT  1.640 0.460 1.960 0.620 ;
        RECT  3.440 0.440 4.260 0.600 ;
        RECT  3.780 0.760 3.940 2.340 ;
        RECT  3.780 1.380 4.080 1.660 ;
        RECT  2.680 2.180 3.600 2.340 ;
        RECT  3.440 0.940 3.600 2.340 ;
        RECT  2.680 0.940 3.600 1.100 ;
        RECT  1.020 2.600 1.960 2.760 ;
        RECT  1.020 2.200 1.180 2.760 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END QDFZRSBHHD

MACRO QDFZSBEHD
    CLASS CORE ;
    FOREIGN QDFZSBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.300 1.420 3.500 1.960 ;
        RECT  3.270 1.480 3.500 1.760 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.420 2.700 1.990 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.500 0.960 10.700 2.120 ;
        RECT  10.480 1.840 10.700 2.120 ;
        RECT  10.480 0.960 10.700 1.240 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.100 1.140 8.300 1.660 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.280 2.800 0.400 ;
        RECT  3.310 -0.280 3.590 0.400 ;
        RECT  6.990 -0.280 7.270 0.400 ;
        RECT  9.850 -0.280 10.130 0.400 ;
        RECT  0.000 -0.280 10.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.470 2.800 3.750 3.480 ;
        RECT  6.980 2.800 7.260 3.480 ;
        RECT  7.740 2.800 8.020 3.480 ;
        RECT  8.980 2.800 9.260 3.480 ;
        RECT  9.900 2.620 10.180 3.480 ;
        RECT  0.000 2.920 10.800 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.480 2.040 9.760 2.320 ;
        RECT  9.480 0.920 9.640 2.320 ;
        RECT  9.240 1.340 10.300 1.620 ;
        RECT  5.210 2.280 5.560 2.440 ;
        RECT  5.210 0.460 5.370 2.440 ;
        RECT  5.850 0.900 7.200 1.060 ;
        RECT  7.040 0.560 7.200 1.060 ;
        RECT  5.850 0.460 6.010 1.060 ;
        RECT  7.040 0.560 7.610 0.720 ;
        RECT  5.210 0.460 6.010 0.620 ;
        RECT  7.450 0.440 9.690 0.600 ;
        RECT  4.890 2.600 5.880 2.760 ;
        RECT  5.720 2.160 5.880 2.760 ;
        RECT  6.980 2.480 9.080 2.640 ;
        RECT  8.920 0.940 9.080 2.640 ;
        RECT  4.890 0.460 5.050 2.760 ;
        RECT  6.980 2.160 7.140 2.640 ;
        RECT  4.510 2.300 5.050 2.460 ;
        RECT  5.720 2.160 7.140 2.320 ;
        RECT  8.920 0.940 9.260 1.100 ;
        RECT  4.730 0.460 5.050 0.680 ;
        RECT  7.300 2.060 8.580 2.220 ;
        RECT  8.300 1.920 8.580 2.220 ;
        RECT  7.300 2.000 7.670 2.220 ;
        RECT  7.510 0.880 7.670 2.220 ;
        RECT  6.510 1.360 7.670 1.520 ;
        RECT  7.360 0.880 7.670 1.520 ;
        RECT  5.530 1.680 5.960 1.980 ;
        RECT  5.530 1.680 7.350 1.840 ;
        RECT  5.530 0.840 5.690 1.980 ;
        RECT  6.170 0.460 6.830 0.740 ;
        RECT  6.040 2.480 6.820 2.760 ;
        RECT  1.480 2.520 2.340 2.680 ;
        RECT  2.180 0.560 2.340 2.680 ;
        RECT  4.570 0.880 4.730 2.040 ;
        RECT  4.410 0.440 4.570 1.040 ;
        RECT  1.600 0.740 2.340 0.900 ;
        RECT  2.180 0.560 3.910 0.720 ;
        RECT  3.750 0.440 4.570 0.600 ;
        RECT  4.090 0.760 4.250 2.400 ;
        RECT  4.090 1.380 4.390 1.660 ;
        RECT  3.030 2.240 3.910 2.460 ;
        RECT  3.750 0.880 3.910 2.460 ;
        RECT  3.090 0.880 3.910 1.160 ;
        RECT  0.900 2.200 2.020 2.360 ;
        RECT  1.860 1.460 2.020 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END QDFZSBEHD

MACRO QDFZSBHHD
    CLASS CORE ;
    FOREIGN QDFZSBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN CK
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.900 1.480 3.260 1.760 ;
        RECT  2.900 1.420 3.100 1.960 ;
        END
    END CK
    PIN TD
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.420 2.700 1.990 ;
        END
    END TD
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.460 1.540 1.740 ;
        RECT  1.300 1.200 1.500 1.790 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 0.800 11.100 2.120 ;
        RECT  10.760 1.840 11.100 2.120 ;
        RECT  10.760 0.800 11.100 1.080 ;
        END
    END Q
    PIN SB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.080 1.380 8.300 1.660 ;
        RECT  8.100 1.140 8.300 1.660 ;
        END
    END SB
    PIN SEL
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.410 0.700 2.240 ;
        RECT  0.420 1.460 0.700 1.740 ;
        END
    END SEL
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 -0.280 2.800 0.400 ;
        RECT  3.190 -0.280 3.470 0.400 ;
        RECT  6.880 -0.280 7.160 0.400 ;
        RECT  8.240 -0.280 8.520 0.400 ;
        RECT  10.140 -0.280 10.420 0.400 ;
        RECT  11.220 -0.280 11.500 0.580 ;
        RECT  0.000 -0.280 11.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.620 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.800 2.800 3.480 ;
        RECT  3.350 2.800 3.630 3.480 ;
        RECT  6.900 2.800 8.480 3.480 ;
        RECT  9.320 2.800 9.600 3.480 ;
        RECT  10.180 2.620 10.460 3.480 ;
        RECT  11.220 2.620 11.500 3.480 ;
        RECT  0.000 2.920 11.600 3.480 ;
        RECT  0.620 2.620 0.900 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  9.620 1.900 10.580 2.060 ;
        RECT  10.420 1.400 10.580 2.060 ;
        RECT  9.620 0.960 9.780 2.060 ;
        RECT  9.460 1.400 9.780 1.680 ;
        RECT  9.560 0.960 9.780 1.680 ;
        RECT  5.090 2.280 5.440 2.440 ;
        RECT  5.090 0.460 5.250 2.440 ;
        RECT  9.940 0.640 10.100 1.620 ;
        RECT  5.730 0.900 7.060 1.060 ;
        RECT  6.900 0.560 7.060 1.060 ;
        RECT  5.730 0.460 5.890 1.060 ;
        RECT  9.640 0.640 10.100 0.800 ;
        RECT  6.900 0.560 9.800 0.720 ;
        RECT  5.090 0.460 5.890 0.620 ;
        RECT  8.760 2.480 9.040 2.760 ;
        RECT  4.770 2.600 5.760 2.760 ;
        RECT  5.600 2.160 5.760 2.760 ;
        RECT  6.880 2.480 9.200 2.640 ;
        RECT  9.040 0.960 9.200 2.640 ;
        RECT  4.770 0.460 4.930 2.760 ;
        RECT  6.880 2.160 7.040 2.640 ;
        RECT  4.390 2.300 4.930 2.460 ;
        RECT  5.600 2.160 7.040 2.320 ;
        RECT  9.040 0.960 9.320 1.240 ;
        RECT  4.610 0.460 4.930 0.680 ;
        RECT  7.200 1.980 7.570 2.280 ;
        RECT  7.410 0.940 7.570 2.280 ;
        RECT  7.200 1.980 8.520 2.140 ;
        RECT  8.200 1.900 8.480 2.140 ;
        RECT  6.410 1.220 6.730 1.480 ;
        RECT  6.410 1.220 7.640 1.380 ;
        RECT  7.360 0.940 7.640 1.380 ;
        RECT  5.410 1.660 5.840 1.980 ;
        RECT  5.410 1.660 7.250 1.820 ;
        RECT  6.970 1.540 7.250 1.820 ;
        RECT  5.410 0.840 5.570 1.980 ;
        RECT  6.140 2.480 6.680 2.760 ;
        RECT  6.070 0.460 6.670 0.740 ;
        RECT  1.480 2.520 2.340 2.680 ;
        RECT  2.180 0.560 2.340 2.680 ;
        RECT  4.450 0.880 4.610 2.040 ;
        RECT  4.290 0.440 4.450 1.040 ;
        RECT  1.600 0.740 2.340 0.900 ;
        RECT  2.180 0.560 3.790 0.720 ;
        RECT  3.630 0.440 4.450 0.600 ;
        RECT  3.970 0.760 4.130 2.450 ;
        RECT  3.970 1.380 4.270 1.660 ;
        RECT  2.870 2.240 3.790 2.400 ;
        RECT  3.630 0.880 3.790 2.400 ;
        RECT  2.870 0.880 3.790 1.040 ;
        RECT  0.900 2.200 2.020 2.360 ;
        RECT  1.860 1.460 2.020 2.360 ;
        RECT  0.100 0.820 0.260 2.320 ;
        RECT  0.100 2.000 0.320 2.280 ;
        RECT  0.900 0.820 1.060 2.360 ;
        RECT  0.100 0.820 1.060 0.980 ;
    END
END QDFZSBHHD

MACRO QDLAHCHD
    CLASS CORE ;
    FOREIGN QDLAHCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.850 5.510 1.130 ;
        RECT  5.300 1.840 5.510 2.120 ;
        RECT  5.300 0.850 5.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.600 ;
        RECT  5.890 -0.280 6.170 0.940 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.850 2.800 6.130 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 0.440 5.030 2.440 ;
        RECT  4.090 0.860 4.250 1.140 ;
        RECT  4.090 0.920 5.030 1.080 ;
        RECT  4.810 0.440 5.090 0.600 ;
        RECT  3.050 2.480 4.630 2.640 ;
        RECT  4.470 1.460 4.630 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.440 3.850 2.320 ;
        RECT  3.690 0.440 3.970 0.600 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  1.290 0.580 2.370 0.740 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  0.100 2.300 2.870 2.460 ;
        RECT  2.710 1.380 2.870 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.330 1.840 2.550 2.120 ;
        RECT  2.390 0.940 2.550 2.120 ;
        RECT  2.330 0.940 2.610 1.100 ;
    END
END QDLAHCHD

MACRO QDLAHEHD
    CLASS CORE ;
    FOREIGN QDLAHEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.300 0.850 5.510 1.130 ;
        RECT  5.300 1.840 5.510 2.120 ;
        RECT  5.300 0.850 5.500 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.980 ;
        RECT  5.890 -0.280 6.170 0.580 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.850 2.800 6.130 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 0.820 5.030 2.440 ;
        RECT  4.030 1.200 4.310 1.420 ;
        RECT  4.030 1.200 5.090 1.360 ;
        RECT  4.810 0.820 5.090 1.360 ;
        RECT  3.050 2.480 4.630 2.640 ;
        RECT  4.470 1.690 4.630 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.820 3.850 2.320 ;
        RECT  3.690 0.820 3.970 0.980 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  1.290 0.580 2.370 0.740 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  0.100 2.300 2.870 2.460 ;
        RECT  2.710 1.380 2.870 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.330 1.850 2.550 2.130 ;
        RECT  2.390 0.940 2.550 2.130 ;
        RECT  2.330 0.940 2.610 1.100 ;
    END
END QDLAHEHD

MACRO QDLAHHHD
    CLASS CORE ;
    FOREIGN QDLAHHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.370 2.150 1.650 ;
        RECT  1.700 1.240 1.900 1.880 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.700 0.850 6.030 1.130 ;
        RECT  5.700 1.840 6.030 2.120 ;
        RECT  5.700 0.850 5.900 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 -0.280 2.050 0.400 ;
        RECT  4.290 -0.280 4.570 0.980 ;
        RECT  5.290 -0.280 5.570 0.580 ;
        RECT  6.330 -0.280 6.610 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.770 2.620 2.050 3.480 ;
        RECT  4.250 2.800 4.530 3.480 ;
        RECT  5.290 2.620 5.570 3.480 ;
        RECT  6.330 2.620 6.610 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.870 0.820 5.030 2.440 ;
        RECT  4.030 1.200 4.310 1.420 ;
        RECT  4.030 1.200 5.090 1.360 ;
        RECT  4.820 0.820 5.090 1.360 ;
        RECT  4.810 0.820 5.090 0.980 ;
        RECT  3.050 2.480 4.700 2.640 ;
        RECT  4.540 1.520 4.700 2.640 ;
        RECT  3.050 0.760 3.210 2.640 ;
        RECT  2.990 0.760 3.210 1.040 ;
        RECT  3.690 2.100 3.970 2.320 ;
        RECT  3.690 0.820 3.850 2.320 ;
        RECT  3.690 0.820 3.970 0.980 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  3.370 0.440 3.530 2.020 ;
        RECT  1.290 0.580 2.370 0.740 ;
        RECT  2.210 0.440 3.530 0.600 ;
        RECT  0.100 2.300 2.890 2.460 ;
        RECT  2.730 1.440 2.890 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 2.220 0.380 2.460 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
        RECT  2.330 1.840 2.550 2.120 ;
        RECT  2.390 0.960 2.550 2.120 ;
    END
END QDLAHHHD

MACRO QDLAHRBCHD
    CLASS CORE ;
    FOREIGN QDLAHRBCHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.340 2.300 1.620 ;
        RECT  2.100 1.000 2.300 1.620 ;
        END
    END RB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.340 2.840 1.620 ;
        RECT  2.500 1.000 2.700 1.620 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.850 6.310 1.130 ;
        RECT  6.100 1.840 6.310 2.120 ;
        RECT  6.100 0.850 6.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.660 ;
        RECT  6.690 -0.280 6.970 0.940 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.490 2.470 2.770 3.480 ;
        RECT  5.220 2.800 5.930 3.480 ;
        RECT  6.650 2.800 6.930 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.670 0.440 5.830 2.410 ;
        RECT  4.890 0.940 5.110 1.220 ;
        RECT  4.890 1.000 5.830 1.160 ;
        RECT  2.930 2.600 5.050 2.760 ;
        RECT  5.270 1.460 5.430 2.640 ;
        RECT  4.890 2.480 5.430 2.640 ;
        RECT  3.890 0.820 4.050 2.760 ;
        RECT  2.930 2.150 3.090 2.760 ;
        RECT  1.930 2.150 2.210 2.370 ;
        RECT  1.930 2.150 3.090 2.310 ;
        RECT  3.710 0.820 4.050 0.980 ;
        RECT  4.530 2.130 4.730 2.410 ;
        RECT  4.530 0.440 4.690 2.410 ;
        RECT  4.530 0.440 4.750 0.720 ;
        RECT  1.290 0.560 1.450 2.120 ;
        RECT  4.210 0.440 4.370 2.060 ;
        RECT  1.290 0.560 2.490 0.720 ;
        RECT  2.330 0.440 4.370 0.600 ;
        RECT  3.270 2.150 3.730 2.310 ;
        RECT  3.570 1.140 3.730 2.310 ;
        RECT  3.350 1.140 3.730 1.300 ;
        RECT  3.350 0.820 3.510 1.300 ;
        RECT  3.230 0.820 3.510 1.040 ;
        RECT  0.100 2.300 0.380 2.520 ;
        RECT  0.100 2.300 1.770 2.460 ;
        RECT  1.610 1.830 1.770 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  1.610 1.830 3.410 1.990 ;
        RECT  3.250 1.510 3.410 1.990 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.660 0.380 0.900 ;
    END
END QDLAHRBCHD

MACRO QDLAHRBEHD
    CLASS CORE ;
    FOREIGN QDLAHRBEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.060 1.340 2.300 1.620 ;
        RECT  2.100 1.000 2.300 1.620 ;
        END
    END RB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.340 2.840 1.620 ;
        RECT  2.500 1.000 2.700 1.620 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.850 6.310 1.130 ;
        RECT  6.100 1.840 6.310 2.120 ;
        RECT  6.100 0.850 6.300 2.120 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.760 ;
        RECT  6.610 -0.280 6.890 0.580 ;
        RECT  0.000 -0.280 7.200 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.490 2.470 2.770 3.480 ;
        RECT  5.220 2.740 5.440 3.480 ;
        RECT  6.650 2.800 6.930 3.480 ;
        RECT  0.000 2.920 7.200 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.670 0.540 5.830 2.450 ;
        RECT  4.890 1.070 5.050 1.350 ;
        RECT  4.890 1.130 5.830 1.290 ;
        RECT  2.930 2.600 5.060 2.760 ;
        RECT  4.900 2.420 5.060 2.760 ;
        RECT  3.890 0.820 4.050 2.760 ;
        RECT  2.930 2.150 3.090 2.760 ;
        RECT  4.900 2.420 5.430 2.580 ;
        RECT  5.270 1.550 5.430 2.580 ;
        RECT  1.930 2.150 2.210 2.370 ;
        RECT  1.930 2.150 3.090 2.310 ;
        RECT  3.710 0.820 4.050 0.980 ;
        RECT  4.530 2.130 4.740 2.410 ;
        RECT  4.530 0.540 4.690 2.410 ;
        RECT  1.290 0.560 1.450 2.120 ;
        RECT  4.210 0.440 4.370 2.060 ;
        RECT  1.290 0.560 2.490 0.720 ;
        RECT  2.330 0.440 4.370 0.600 ;
        RECT  3.270 2.150 3.730 2.310 ;
        RECT  3.570 1.140 3.730 2.310 ;
        RECT  3.350 1.140 3.730 1.300 ;
        RECT  3.350 0.820 3.510 1.300 ;
        RECT  3.230 0.820 3.510 1.040 ;
        RECT  0.100 2.300 1.770 2.460 ;
        RECT  1.610 1.830 1.770 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  1.610 1.830 3.410 1.990 ;
        RECT  3.250 1.510 3.410 1.990 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END QDLAHRBEHD

MACRO QDLAHRBHHD
    CLASS CORE ;
    FOREIGN QDLAHRBHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN RB
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.100 1.000 2.300 1.650 ;
        END
    END RB
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.370 2.970 1.650 ;
        RECT  2.500 1.000 2.700 1.650 ;
        END
    END D
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.900 0.900 7.100 2.300 ;
        RECT  6.700 2.100 7.100 2.300 ;
        RECT  6.660 0.900 7.100 1.100 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.890 -0.280 2.170 0.400 ;
        RECT  5.090 -0.280 5.370 0.980 ;
        RECT  6.140 -0.280 6.420 0.580 ;
        RECT  7.180 -0.280 7.460 0.580 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.520 2.620 2.800 3.480 ;
        RECT  5.240 2.320 5.460 3.480 ;
        RECT  6.180 2.620 6.460 3.480 ;
        RECT  7.220 2.620 7.500 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.760 0.820 5.920 2.400 ;
        RECT  4.890 1.140 5.110 1.420 ;
        RECT  4.890 1.200 5.920 1.360 ;
        RECT  5.660 0.820 5.940 0.980 ;
        RECT  2.970 2.570 5.080 2.730 ;
        RECT  4.920 1.940 5.080 2.730 ;
        RECT  3.930 0.760 4.090 2.730 ;
        RECT  2.970 2.300 3.130 2.730 ;
        RECT  1.930 2.300 3.130 2.460 ;
        RECT  4.920 1.940 5.590 2.100 ;
        RECT  5.370 1.560 5.590 2.100 ;
        RECT  4.570 2.130 4.760 2.410 ;
        RECT  4.570 0.760 4.730 2.410 ;
        RECT  1.290 0.580 1.450 2.120 ;
        RECT  4.250 0.440 4.410 2.070 ;
        RECT  1.290 0.580 2.490 0.740 ;
        RECT  2.330 0.440 4.410 0.600 ;
        RECT  3.310 2.240 3.770 2.400 ;
        RECT  3.610 0.940 3.770 2.400 ;
        RECT  3.190 0.940 3.770 1.100 ;
        RECT  3.190 0.820 3.410 1.100 ;
        RECT  0.100 2.300 1.770 2.460 ;
        RECT  1.610 1.920 1.770 2.460 ;
        RECT  0.850 0.740 1.010 2.460 ;
        RECT  0.100 2.220 0.380 2.460 ;
        RECT  1.610 1.920 3.450 2.080 ;
        RECT  3.290 1.480 3.450 2.080 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END QDLAHRBHHD

MACRO QDLAHSEHD
    CLASS CORE ;
    FOREIGN QDLAHSEHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.460 2.710 1.740 ;
        RECT  2.500 1.460 2.700 2.020 ;
        END
    END D
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 2.000 1.740 ;
        RECT  1.700 1.400 1.900 2.020 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  6.100 0.850 6.300 2.120 ;
        RECT  5.940 1.840 6.300 2.120 ;
        RECT  5.940 0.850 6.300 1.130 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.280 2.060 0.460 ;
        RECT  4.880 -0.280 5.160 0.760 ;
        RECT  6.400 -0.280 6.680 0.580 ;
        RECT  0.000 -0.280 6.800 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.710 2.620 1.990 3.480 ;
        RECT  5.010 2.740 5.230 3.480 ;
        RECT  6.400 2.620 6.680 3.480 ;
        RECT  0.000 2.920 6.800 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.460 0.540 5.620 2.450 ;
        RECT  4.680 1.070 4.840 1.350 ;
        RECT  4.680 1.130 5.620 1.290 ;
        RECT  3.680 2.600 4.850 2.760 ;
        RECT  4.690 2.420 4.850 2.760 ;
        RECT  3.680 0.760 3.840 2.760 ;
        RECT  4.690 2.420 5.220 2.580 ;
        RECT  5.060 1.550 5.220 2.580 ;
        RECT  1.710 0.950 2.750 1.110 ;
        RECT  2.590 0.760 2.750 1.110 ;
        RECT  3.540 0.760 3.840 0.980 ;
        RECT  2.590 0.760 3.840 0.920 ;
        RECT  4.320 2.130 4.530 2.410 ;
        RECT  4.320 0.540 4.480 2.410 ;
        RECT  1.290 0.630 1.450 2.120 ;
        RECT  4.000 0.440 4.160 2.060 ;
        RECT  1.290 0.630 2.410 0.790 ;
        RECT  2.250 0.440 2.410 0.790 ;
        RECT  2.250 0.440 4.160 0.600 ;
        RECT  2.980 2.600 3.520 2.760 ;
        RECT  3.360 1.140 3.520 2.760 ;
        RECT  2.980 1.140 3.520 1.300 ;
        RECT  2.980 1.080 3.260 1.300 ;
        RECT  0.100 2.280 3.200 2.440 ;
        RECT  3.040 1.510 3.200 2.440 ;
        RECT  0.850 0.740 1.010 2.440 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END QDLAHSEHD

MACRO QDLAHSHHD
    CLASS CORE ;
    FOREIGN QDLAHSHHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN G
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.370 0.420 1.650 ;
        RECT  0.100 1.240 0.300 1.880 ;
        END
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.500 1.460 2.710 1.740 ;
        RECT  2.500 1.460 2.700 2.020 ;
        END
    END D
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.460 2.000 1.740 ;
        RECT  1.700 1.400 1.900 2.020 ;
        END
    END S
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.940 0.920 7.300 1.080 ;
        RECT  5.940 2.120 7.300 2.280 ;
        RECT  6.500 0.920 6.700 2.280 ;
        END
    END Q
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.840 -0.280 2.060 0.460 ;
        RECT  4.940 -0.280 5.220 0.760 ;
        RECT  6.460 -0.280 6.740 0.580 ;
        RECT  0.000 -0.280 7.600 0.280 ;
        RECT  0.660 -0.280 0.940 0.580 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.710 2.620 1.990 3.480 ;
        RECT  4.960 2.740 5.180 3.480 ;
        RECT  6.460 2.620 6.740 3.480 ;
        RECT  0.000 2.920 7.600 3.480 ;
        RECT  0.660 2.620 0.940 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.520 0.540 5.680 2.450 ;
        RECT  4.680 1.070 4.840 1.350 ;
        RECT  4.680 1.130 5.680 1.290 ;
        RECT  3.680 2.600 4.800 2.760 ;
        RECT  4.640 2.420 4.800 2.760 ;
        RECT  3.680 0.760 3.840 2.760 ;
        RECT  4.640 2.420 5.280 2.580 ;
        RECT  5.120 1.550 5.280 2.580 ;
        RECT  1.710 0.950 2.750 1.110 ;
        RECT  2.590 0.760 2.750 1.110 ;
        RECT  3.540 0.760 3.840 0.980 ;
        RECT  2.590 0.760 3.840 0.920 ;
        RECT  4.260 2.190 4.480 2.440 ;
        RECT  4.360 0.540 4.520 2.310 ;
        RECT  4.320 2.130 4.520 2.310 ;
        RECT  4.320 0.540 4.520 0.820 ;
        RECT  1.290 0.630 1.450 2.120 ;
        RECT  4.000 0.440 4.160 2.060 ;
        RECT  4.000 1.740 4.200 2.020 ;
        RECT  1.290 0.630 2.410 0.790 ;
        RECT  2.250 0.440 2.410 0.790 ;
        RECT  2.250 0.440 4.160 0.600 ;
        RECT  2.980 2.600 3.520 2.760 ;
        RECT  3.360 1.140 3.520 2.760 ;
        RECT  2.980 1.140 3.520 1.300 ;
        RECT  2.980 1.080 3.260 1.300 ;
        RECT  0.100 2.280 3.200 2.440 ;
        RECT  3.040 1.510 3.200 2.440 ;
        RECT  0.850 0.740 1.010 2.440 ;
        RECT  0.100 0.740 1.010 0.900 ;
        RECT  0.100 0.720 0.380 0.900 ;
    END
END QDLAHSHHD

MACRO TIE0DHD
    CLASS CORE ;
    FOREIGN TIE0DHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.340 0.570 0.540 1.210 ;
        RECT  0.100 0.900 0.540 1.210 ;
        RECT  0.100 0.900 0.300 1.960 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        RECT  0.820 -0.280 1.100 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        RECT  0.820 2.010 1.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.360 2.200 0.660 2.480 ;
        RECT  0.500 1.460 0.660 2.480 ;
    END
END TIE0DHD

MACRO TIE0HHD
    CLASS CORE ;
    FOREIGN TIE0HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.660 0.900 1.500 1.100 ;
        RECT  1.300 0.900 1.500 1.960 ;
        RECT  0.660 0.600 0.860 1.240 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.700 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 0.380 1.240 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.200 1.420 3.480 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 1.900 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.680 1.460 0.840 2.540 ;
    END
END TIE0HHD

MACRO TIE0KHD
    CLASS CORE ;
    FOREIGN TIE0KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 0.600 1.900 1.320 ;
        RECT  0.660 1.120 2.700 1.320 ;
        RECT  2.500 1.120 2.700 2.360 ;
        RECT  0.660 0.600 0.860 1.320 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.900 ;
        RECT  2.180 -0.280 2.460 0.900 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.100 -0.280 0.380 1.240 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 1.980 1.420 3.480 ;
        RECT  2.180 2.560 2.460 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 1.900 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.720 1.520 1.880 2.640 ;
        RECT  0.680 1.520 0.840 2.540 ;
        RECT  0.680 1.520 1.880 1.680 ;
    END
END TIE0KHD

MACRO TIE1DHD
    CLASS CORE ;
    FOREIGN TIE1DHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 2.020 0.540 2.300 ;
        RECT  0.340 2.020 0.540 2.660 ;
        RECT  0.100 1.240 0.300 2.300 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.280 1.200 0.280 ;
        RECT  0.820 -0.280 1.100 1.210 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 2.920 1.200 3.480 ;
        RECT  0.820 2.010 1.100 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.500 0.740 0.660 1.620 ;
        RECT  0.360 0.740 0.660 1.020 ;
    END
END TIE1DHD

MACRO TIE1HHD
    CLASS CORE ;
    FOREIGN TIE1HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.600 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 0.840 1.500 1.980 ;
        RECT  0.660 1.780 1.500 1.980 ;
        RECT  0.660 1.780 0.860 2.540 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 0.640 ;
        RECT  0.000 -0.280 1.600 0.280 ;
        RECT  0.100 -0.280 0.380 1.240 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.200 1.420 3.480 ;
        RECT  0.000 2.920 1.600 3.480 ;
        RECT  0.100 1.900 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.680 0.600 0.840 1.620 ;
    END
END TIE1HHD

MACRO TIE1KHD
    CLASS CORE ;
    FOREIGN TIE1KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.700 1.720 1.900 2.640 ;
        RECT  2.500 0.840 2.700 1.920 ;
        RECT  0.660 1.720 2.700 1.920 ;
        RECT  0.660 1.720 0.860 2.540 ;
        END
    END O
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 -0.280 1.420 1.110 ;
        RECT  2.180 -0.280 2.460 0.640 ;
        RECT  0.000 -0.280 2.800 0.280 ;
        RECT  0.100 -0.280 0.380 1.240 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.140 2.080 1.420 3.480 ;
        RECT  2.180 2.100 2.460 3.480 ;
        RECT  0.000 2.920 2.800 3.480 ;
        RECT  0.100 1.900 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.680 1.400 1.880 1.560 ;
        RECT  1.720 0.500 1.880 1.560 ;
        RECT  0.680 0.500 0.840 1.560 ;
    END
END TIE1KHD

MACRO XNR2CHD
    CLASS CORE ;
    FOREIGN XNR2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 2.140 4.300 2.420 ;
        RECT  4.100 0.440 4.300 2.680 ;
        RECT  4.080 0.600 4.300 0.880 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.640 0.700 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.860 0.800 1.140 1.080 ;
        RECT  3.450 -0.280 3.730 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.920 -0.280 1.080 1.080 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.450 2.800 3.730 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.600 3.240 2.760 ;
        RECT  3.720 0.560 3.880 2.640 ;
        RECT  3.080 2.480 3.880 2.640 ;
        RECT  2.080 2.100 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 3.880 0.720 ;
        RECT  2.620 2.120 2.900 2.320 ;
        RECT  2.620 2.120 3.560 2.280 ;
        RECT  3.400 0.880 3.560 2.280 ;
        RECT  2.880 0.880 3.560 1.040 ;
        RECT  1.440 1.320 1.600 2.420 ;
        RECT  1.440 1.320 3.240 1.480 ;
        RECT  2.980 1.200 3.240 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.730 1.920 2.760 ;
        RECT  0.120 2.480 1.280 2.640 ;
        RECT  0.120 2.280 0.340 2.640 ;
        RECT  0.120 0.520 0.280 2.640 ;
        RECT  2.700 1.680 2.980 1.960 ;
        RECT  1.760 1.730 2.980 1.890 ;
        RECT  0.120 0.800 0.340 1.080 ;
    END
END XNR2CHD

MACRO XNR2EHD
    CLASS CORE ;
    FOREIGN XNR2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 2.420 4.300 2.700 ;
        RECT  4.100 0.440 4.300 2.740 ;
        RECT  4.080 0.480 4.300 0.760 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.640 0.700 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.860 0.800 1.140 1.080 ;
        RECT  3.450 -0.280 3.730 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.920 -0.280 1.080 1.080 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.450 2.800 3.730 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.600 3.240 2.760 ;
        RECT  3.720 0.560 3.880 2.640 ;
        RECT  3.080 2.480 3.880 2.640 ;
        RECT  2.080 2.140 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 3.880 0.720 ;
        RECT  2.620 2.120 2.900 2.360 ;
        RECT  2.620 2.120 3.560 2.280 ;
        RECT  3.400 0.880 3.560 2.280 ;
        RECT  2.880 0.880 3.560 1.040 ;
        RECT  1.440 1.320 1.600 2.420 ;
        RECT  1.430 1.320 3.240 1.480 ;
        RECT  2.980 1.200 3.240 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.760 1.920 2.760 ;
        RECT  0.120 2.480 1.280 2.640 ;
        RECT  0.120 2.320 0.340 2.640 ;
        RECT  0.120 0.520 0.280 2.640 ;
        RECT  1.760 1.760 2.980 1.920 ;
        RECT  0.120 0.800 0.340 1.080 ;
    END
END XNR2EHD

MACRO XNR2HHD
    CLASS CORE ;
    FOREIGN XNR2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.500 4.700 2.700 ;
        RECT  4.260 2.500 4.700 2.700 ;
        RECT  4.260 0.500 4.700 0.700 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.640 0.700 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.630 -0.280 3.910 0.400 ;
        RECT  4.880 -0.280 5.040 0.500 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.920 -0.280 1.080 1.040 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.630 2.800 3.910 3.480 ;
        RECT  4.880 2.700 5.040 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.600 3.420 2.760 ;
        RECT  3.900 0.560 4.060 2.640 ;
        RECT  3.260 2.480 4.060 2.640 ;
        RECT  2.080 2.140 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 4.060 0.720 ;
        RECT  2.620 2.120 2.900 2.360 ;
        RECT  2.620 2.120 3.740 2.280 ;
        RECT  3.580 0.880 3.740 2.280 ;
        RECT  2.880 0.880 3.740 1.040 ;
        RECT  1.440 1.320 1.600 2.420 ;
        RECT  1.440 1.320 3.420 1.480 ;
        RECT  3.160 1.200 3.420 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.660 1.920 2.760 ;
        RECT  0.120 2.480 1.280 2.640 ;
        RECT  0.120 2.320 0.340 2.640 ;
        RECT  0.120 0.520 0.280 2.640 ;
        RECT  1.760 1.660 2.980 1.820 ;
        RECT  0.120 0.800 0.340 1.080 ;
    END
END XNR2HHD

MACRO XNR2KHD
    CLASS CORE ;
    FOREIGN XNR2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.560 0.460 5.900 0.740 ;
        RECT  4.500 1.700 5.900 1.900 ;
        RECT  5.700 0.460 5.900 2.740 ;
        RECT  5.560 2.460 5.900 2.740 ;
        RECT  4.500 0.460 4.700 2.740 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 0.600 1.360 0.760 ;
        RECT  1.200 0.520 2.300 0.680 ;
        RECT  2.020 0.440 2.300 0.680 ;
        RECT  0.500 0.600 0.700 1.560 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.340 1.180 1.620 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.890 -0.280 4.170 0.400 ;
        RECT  5.040 -0.280 5.200 0.640 ;
        RECT  6.080 -0.280 6.240 0.680 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.750 -0.280 1.030 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.890 2.800 4.170 3.480 ;
        RECT  5.040 2.560 5.200 3.480 ;
        RECT  6.080 2.520 6.240 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.480 4.320 2.640 ;
        RECT  4.160 0.560 4.320 2.640 ;
        RECT  2.080 2.140 2.240 2.640 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 4.320 0.720 ;
        RECT  2.620 2.120 4.000 2.280 ;
        RECT  3.840 0.880 4.000 2.280 ;
        RECT  2.840 0.880 4.000 1.040 ;
        RECT  1.440 1.240 1.600 2.220 ;
        RECT  3.420 1.240 3.680 1.640 ;
        RECT  1.440 1.240 3.680 1.400 ;
        RECT  1.860 0.960 2.020 1.400 ;
        RECT  0.120 2.480 1.920 2.640 ;
        RECT  1.760 1.560 1.920 2.640 ;
        RECT  0.120 2.320 0.340 2.640 ;
        RECT  0.120 0.460 0.280 2.640 ;
        RECT  1.760 1.560 1.960 1.840 ;
        RECT  1.760 1.560 2.980 1.720 ;
        RECT  0.120 0.460 0.340 0.740 ;
    END
END XNR2KHD

MACRO XNR3CHD
    CLASS CORE ;
    FOREIGN XNR3CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.440 0.710 8.600 0.990 ;
        RECT  8.500 0.720 8.700 2.530 ;
        RECT  8.440 2.240 8.700 2.520 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.640 0.420 1.920 ;
        RECT  0.100 1.640 0.300 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.640 7.900 2.280 ;
        RECT  7.660 1.830 7.900 2.110 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.620 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  7.820 2.800 8.100 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 0.440 6.480 2.300 ;
        RECT  8.080 0.560 8.240 1.620 ;
        RECT  7.320 0.560 8.240 0.720 ;
        RECT  6.320 0.440 7.480 0.600 ;
        RECT  7.320 0.960 7.480 2.720 ;
        RECT  7.180 1.440 7.480 1.720 ;
        RECT  5.480 2.600 7.000 2.760 ;
        RECT  6.840 0.780 7.000 2.760 ;
        RECT  5.480 0.760 5.640 2.760 ;
        RECT  4.600 0.760 4.760 2.300 ;
        RECT  4.600 0.760 5.640 0.920 ;
        RECT  5.800 0.440 5.960 2.300 ;
        RECT  3.520 0.440 3.680 2.120 ;
        RECT  3.520 0.440 5.960 0.600 ;
        RECT  2.880 2.600 5.320 2.760 ;
        RECT  5.160 1.080 5.320 2.760 ;
        RECT  2.880 0.840 3.040 2.760 ;
        RECT  3.200 2.280 4.240 2.440 ;
        RECT  4.080 0.780 4.240 2.440 ;
        RECT  1.140 2.160 2.280 2.320 ;
        RECT  3.200 0.440 3.360 2.440 ;
        RECT  2.120 0.780 2.280 2.320 ;
        RECT  1.100 0.780 2.300 0.940 ;
        RECT  2.140 0.440 2.300 0.940 ;
        RECT  2.140 0.440 3.360 0.600 ;
        RECT  0.720 2.480 2.720 2.640 ;
        RECT  2.460 2.360 2.720 2.640 ;
        RECT  0.720 0.920 0.880 2.640 ;
    END
END XNR3CHD

MACRO XNR3EHD
    CLASS CORE ;
    FOREIGN XNR3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.480 0.710 8.700 2.280 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.420 1.620 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.320 7.900 1.960 ;
        RECT  7.660 1.340 7.900 1.620 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.620 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  7.820 2.800 8.100 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 0.440 6.480 2.300 ;
        RECT  8.140 0.560 8.300 1.660 ;
        RECT  7.320 0.560 8.300 0.720 ;
        RECT  6.320 0.440 7.480 0.600 ;
        RECT  7.320 0.960 7.480 2.720 ;
        RECT  7.180 1.440 7.480 1.720 ;
        RECT  5.480 2.600 7.000 2.760 ;
        RECT  6.840 0.780 7.000 2.760 ;
        RECT  5.480 0.760 5.640 2.760 ;
        RECT  4.600 0.760 4.760 2.300 ;
        RECT  4.600 0.760 5.640 0.920 ;
        RECT  5.800 0.440 5.960 2.300 ;
        RECT  3.520 0.440 3.680 2.120 ;
        RECT  3.520 0.440 5.960 0.600 ;
        RECT  2.880 2.600 5.320 2.760 ;
        RECT  5.160 1.080 5.320 2.760 ;
        RECT  2.880 0.760 3.040 2.760 ;
        RECT  2.800 0.760 3.040 1.040 ;
        RECT  3.200 2.280 4.240 2.440 ;
        RECT  4.080 0.780 4.240 2.440 ;
        RECT  1.140 2.160 2.300 2.320 ;
        RECT  2.140 0.440 2.300 2.320 ;
        RECT  3.200 0.440 3.360 2.440 ;
        RECT  1.100 0.780 2.300 0.940 ;
        RECT  2.140 0.440 3.360 0.600 ;
        RECT  0.720 2.480 2.720 2.640 ;
        RECT  2.460 2.360 2.720 2.640 ;
        RECT  0.720 0.920 0.880 2.640 ;
    END
END XNR3EHD

MACRO XNR4EHD
    CLASS CORE ;
    FOREIGN XNR4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 0.900 7.900 2.700 ;
        RECT  7.500 2.500 7.900 2.700 ;
        RECT  7.500 0.900 7.900 1.100 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 1.640 11.500 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.240 11.100 1.880 ;
        RECT  10.820 1.240 11.100 1.520 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.640 0.700 2.280 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.510 -0.280 3.790 0.400 ;
        RECT  6.890 -0.280 7.170 0.400 ;
        RECT  8.210 -0.280 8.490 0.400 ;
        RECT  10.920 -0.280 11.080 1.080 ;
        RECT  10.860 0.800 11.140 1.080 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.860 -0.280 1.140 1.020 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.510 2.800 3.790 3.480 ;
        RECT  6.880 2.800 7.160 3.480 ;
        RECT  8.210 2.800 8.490 3.480 ;
        RECT  11.040 2.800 11.320 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.080 2.600 10.880 2.760 ;
        RECT  11.720 0.800 11.880 2.640 ;
        RECT  10.720 2.480 11.880 2.640 ;
        RECT  11.660 2.320 11.880 2.640 ;
        RECT  10.080 1.720 10.240 2.760 ;
        RECT  9.020 1.720 9.300 1.940 ;
        RECT  9.020 1.720 10.240 1.880 ;
        RECT  11.660 0.800 11.880 1.080 ;
        RECT  10.400 1.320 10.560 2.360 ;
        RECT  8.720 1.320 10.570 1.480 ;
        RECT  10.120 0.780 10.280 1.480 ;
        RECT  8.720 1.200 8.980 1.480 ;
        RECT  8.760 2.600 9.920 2.760 ;
        RECT  9.760 2.140 9.920 2.760 ;
        RECT  8.060 2.480 8.920 2.640 ;
        RECT  8.060 0.560 8.220 2.640 ;
        RECT  9.360 0.880 9.640 1.040 ;
        RECT  9.360 0.560 9.520 1.040 ;
        RECT  6.450 0.560 9.520 0.720 ;
        RECT  6.450 0.480 6.730 0.720 ;
        RECT  9.100 2.120 9.380 2.360 ;
        RECT  8.380 2.120 9.380 2.280 ;
        RECT  8.380 0.880 8.540 2.280 ;
        RECT  8.380 0.880 9.120 1.040 ;
        RECT  4.450 2.600 6.670 2.760 ;
        RECT  7.150 1.400 7.310 2.640 ;
        RECT  6.510 2.480 7.310 2.640 ;
        RECT  5.410 2.100 5.570 2.760 ;
        RECT  4.450 0.920 4.610 2.760 ;
        RECT  4.450 0.920 4.890 1.080 ;
        RECT  4.730 0.440 4.890 1.080 ;
        RECT  5.430 0.880 5.970 1.040 ;
        RECT  5.430 0.440 5.590 1.040 ;
        RECT  4.730 0.440 5.590 0.600 ;
        RECT  5.950 2.120 6.230 2.320 ;
        RECT  5.950 2.120 6.990 2.280 ;
        RECT  6.830 0.880 6.990 2.280 ;
        RECT  6.210 0.880 6.990 1.040 ;
        RECT  4.770 1.320 4.930 2.420 ;
        RECT  4.770 1.320 6.670 1.480 ;
        RECT  6.410 1.200 6.670 1.480 ;
        RECT  5.050 0.780 5.210 1.480 ;
        RECT  5.170 1.760 6.310 1.920 ;
        RECT  4.130 0.440 4.290 2.680 ;
        RECT  4.130 0.440 4.490 0.600 ;
        RECT  2.080 2.600 3.240 2.760 ;
        RECT  3.790 0.560 3.950 2.640 ;
        RECT  3.080 2.480 3.950 2.640 ;
        RECT  2.080 2.140 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 3.950 0.720 ;
        RECT  2.620 2.120 2.900 2.360 ;
        RECT  2.620 2.120 3.620 2.280 ;
        RECT  3.460 0.880 3.620 2.280 ;
        RECT  2.880 0.880 3.620 1.040 ;
        RECT  1.440 1.320 1.600 2.360 ;
        RECT  1.430 1.320 3.280 1.480 ;
        RECT  3.000 1.200 3.280 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.720 1.920 2.760 ;
        RECT  0.120 2.480 1.280 2.640 ;
        RECT  0.120 2.320 0.340 2.640 ;
        RECT  0.120 0.800 0.280 2.640 ;
        RECT  2.700 1.720 2.980 1.940 ;
        RECT  1.760 1.720 2.980 1.880 ;
        RECT  0.120 0.800 0.340 1.080 ;
    END
END XNR4EHD

MACRO XOR2CHD
    CLASS CORE ;
    FOREIGN XOR2CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 2.140 4.300 2.420 ;
        RECT  4.100 0.440 4.300 2.680 ;
        RECT  4.080 0.600 4.300 0.880 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 2.480 1.280 2.640 ;
        RECT  1.760 1.730 1.920 2.760 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.730 2.980 1.890 ;
        RECT  2.700 1.680 2.980 1.960 ;
        RECT  0.500 1.640 0.700 2.640 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.860 0.800 1.140 1.080 ;
        RECT  3.450 -0.280 3.730 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.920 -0.280 1.080 1.080 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.450 2.800 3.730 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.600 3.240 2.760 ;
        RECT  3.720 0.560 3.880 2.640 ;
        RECT  3.080 2.480 3.880 2.640 ;
        RECT  2.080 2.100 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 3.880 0.720 ;
        RECT  2.620 2.120 2.900 2.320 ;
        RECT  2.620 2.120 3.560 2.280 ;
        RECT  3.400 0.880 3.560 2.280 ;
        RECT  2.880 0.880 3.560 1.040 ;
        RECT  1.440 1.320 1.600 2.420 ;
        RECT  1.440 1.320 3.240 1.480 ;
        RECT  2.980 1.200 3.240 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  0.120 0.480 0.280 2.540 ;
        RECT  0.120 2.220 0.340 2.500 ;
        RECT  0.120 0.480 0.340 1.080 ;
        RECT  0.120 0.480 0.400 0.640 ;
    END
END XOR2CHD

MACRO XOR2EHD
    CLASS CORE ;
    FOREIGN XOR2EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.080 2.420 4.300 2.700 ;
        RECT  4.100 0.440 4.300 2.740 ;
        RECT  4.080 0.480 4.300 0.760 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 2.480 1.280 2.640 ;
        RECT  1.760 1.740 1.920 2.760 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.740 2.980 1.900 ;
        RECT  0.500 1.640 0.700 2.640 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.860 0.800 1.140 1.080 ;
        RECT  3.450 -0.280 3.730 0.400 ;
        RECT  0.000 -0.280 4.400 0.280 ;
        RECT  0.920 -0.280 1.080 1.080 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.450 2.800 3.730 3.480 ;
        RECT  0.000 2.920 4.400 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.600 3.240 2.760 ;
        RECT  3.720 0.560 3.880 2.640 ;
        RECT  3.080 2.480 3.880 2.640 ;
        RECT  2.080 2.140 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 3.880 0.720 ;
        RECT  2.620 2.120 2.900 2.360 ;
        RECT  2.620 2.120 3.560 2.280 ;
        RECT  3.400 0.880 3.560 2.280 ;
        RECT  2.880 0.880 3.560 1.040 ;
        RECT  1.440 1.320 1.600 2.380 ;
        RECT  1.430 1.320 3.240 1.480 ;
        RECT  2.980 1.200 3.240 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  0.120 2.320 0.340 2.600 ;
        RECT  0.120 0.480 0.280 2.600 ;
        RECT  0.120 0.480 0.340 1.080 ;
        RECT  0.120 0.480 0.400 0.640 ;
    END
END XOR2EHD

MACRO XOR2HHD
    CLASS CORE ;
    FOREIGN XOR2HHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.200 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.500 0.500 4.700 2.700 ;
        RECT  4.260 2.500 4.700 2.700 ;
        RECT  4.260 0.500 4.700 0.700 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 2.480 1.280 2.640 ;
        RECT  1.760 1.660 1.920 2.760 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.660 2.980 1.820 ;
        RECT  0.500 1.640 0.700 2.640 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.630 -0.280 3.910 0.400 ;
        RECT  4.880 -0.280 5.040 0.500 ;
        RECT  0.000 -0.280 5.200 0.280 ;
        RECT  0.820 -0.280 1.100 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.630 2.800 3.910 3.480 ;
        RECT  4.880 2.700 5.040 3.480 ;
        RECT  0.000 2.920 5.200 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.600 3.420 2.760 ;
        RECT  3.900 0.560 4.060 2.640 ;
        RECT  3.260 2.480 4.060 2.640 ;
        RECT  2.080 2.140 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 4.060 0.720 ;
        RECT  2.620 2.120 2.900 2.360 ;
        RECT  2.620 2.120 3.740 2.280 ;
        RECT  3.580 0.880 3.740 2.280 ;
        RECT  2.880 0.880 3.740 1.040 ;
        RECT  1.440 1.320 1.600 2.370 ;
        RECT  1.440 1.320 3.420 1.480 ;
        RECT  3.160 1.200 3.420 1.480 ;
        RECT  1.720 0.780 1.880 1.480 ;
        RECT  0.120 2.450 0.340 2.730 ;
        RECT  0.120 0.560 0.280 2.730 ;
        RECT  0.120 0.560 0.340 0.980 ;
        RECT  0.120 0.560 1.480 0.720 ;
        RECT  1.320 0.440 2.120 0.600 ;
    END
END XOR2HHD

MACRO XOR2KHD
    CLASS CORE ;
    FOREIGN XOR2KHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.400 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.560 0.460 5.900 0.740 ;
        RECT  4.500 1.700 5.900 1.900 ;
        RECT  5.700 0.460 5.900 2.740 ;
        RECT  5.560 2.460 5.900 2.740 ;
        RECT  4.500 0.460 4.700 2.740 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.760 1.560 1.920 2.640 ;
        RECT  0.500 2.480 1.920 2.640 ;
        RECT  1.760 1.560 1.980 1.840 ;
        RECT  1.760 1.620 2.980 1.780 ;
        RECT  0.500 1.280 0.700 2.640 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.280 1.180 1.560 ;
        RECT  0.900 0.920 1.100 1.560 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.890 -0.280 4.170 0.400 ;
        RECT  5.040 -0.280 5.200 0.640 ;
        RECT  6.080 -0.280 6.240 0.680 ;
        RECT  0.000 -0.280 6.400 0.280 ;
        RECT  0.750 -0.280 1.030 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.890 2.800 4.170 3.480 ;
        RECT  5.040 2.560 5.200 3.480 ;
        RECT  6.080 2.520 6.240 3.480 ;
        RECT  0.000 2.920 6.400 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.080 2.480 4.320 2.640 ;
        RECT  4.160 0.560 4.320 2.640 ;
        RECT  2.080 2.140 2.240 2.640 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 4.320 0.720 ;
        RECT  2.620 2.120 4.000 2.280 ;
        RECT  3.840 0.880 4.000 2.280 ;
        RECT  2.840 0.880 4.000 1.040 ;
        RECT  1.440 1.240 1.600 2.220 ;
        RECT  3.380 1.240 3.660 1.540 ;
        RECT  1.440 1.240 3.660 1.400 ;
        RECT  1.860 0.880 2.020 1.400 ;
        RECT  0.120 2.000 0.340 2.280 ;
        RECT  0.120 0.560 0.280 2.280 ;
        RECT  0.120 0.560 0.340 1.040 ;
        RECT  0.120 0.560 1.480 0.720 ;
        RECT  2.020 0.440 2.300 0.680 ;
        RECT  1.320 0.520 2.300 0.680 ;
    END
END XOR2KHD

MACRO XOR3CHD
    CLASS CORE ;
    FOREIGN XOR3CHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.480 0.920 8.700 2.680 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.640 0.420 1.920 ;
        RECT  0.100 1.640 0.300 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.640 7.900 2.280 ;
        RECT  7.660 1.830 7.900 2.110 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.620 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  7.820 2.800 8.100 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 0.440 6.480 2.300 ;
        RECT  8.080 0.560 8.240 1.660 ;
        RECT  7.320 0.560 8.240 0.720 ;
        RECT  6.320 0.440 7.480 0.600 ;
        RECT  7.320 0.960 7.480 2.720 ;
        RECT  7.180 1.440 7.480 1.720 ;
        RECT  5.480 2.600 7.000 2.760 ;
        RECT  6.840 0.780 7.000 2.760 ;
        RECT  5.480 0.760 5.640 2.760 ;
        RECT  4.600 0.760 4.760 2.300 ;
        RECT  4.600 0.760 5.640 0.920 ;
        RECT  5.800 0.440 5.960 2.300 ;
        RECT  3.520 0.440 3.680 2.120 ;
        RECT  3.520 0.440 5.960 0.600 ;
        RECT  2.880 2.600 5.320 2.760 ;
        RECT  5.160 1.080 5.320 2.760 ;
        RECT  2.880 0.760 3.040 2.760 ;
        RECT  2.800 0.760 3.040 1.040 ;
        RECT  3.200 2.280 4.240 2.440 ;
        RECT  4.080 0.780 4.240 2.440 ;
        RECT  1.140 2.160 2.300 2.320 ;
        RECT  2.140 0.440 2.300 2.320 ;
        RECT  3.200 0.440 3.360 2.440 ;
        RECT  1.100 0.780 2.300 0.940 ;
        RECT  2.140 0.440 3.360 0.600 ;
        RECT  0.720 2.480 2.720 2.640 ;
        RECT  2.460 2.360 2.720 2.640 ;
        RECT  0.720 0.920 0.880 2.640 ;
    END
END XOR3CHD

MACRO XOR3EHD
    CLASS CORE ;
    FOREIGN XOR3EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.800 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  8.480 0.460 8.700 2.740 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.100 1.340 0.420 1.620 ;
        RECT  0.100 1.320 0.300 1.880 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.300 1.240 1.500 1.880 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 1.320 7.900 1.960 ;
        RECT  7.660 1.340 7.900 1.620 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 -0.280 1.980 0.620 ;
        RECT  7.820 -0.280 8.100 0.400 ;
        RECT  0.000 -0.280 8.800 0.280 ;
        RECT  0.100 -0.280 0.380 0.400 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.700 2.800 1.980 3.480 ;
        RECT  7.820 2.800 8.100 3.480 ;
        RECT  0.000 2.920 8.800 3.480 ;
        RECT  0.100 2.800 0.380 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  6.320 0.440 6.480 2.300 ;
        RECT  8.140 0.560 8.300 1.660 ;
        RECT  7.320 0.560 8.300 0.720 ;
        RECT  6.320 0.440 7.480 0.600 ;
        RECT  7.320 0.960 7.480 2.720 ;
        RECT  7.180 1.440 7.480 1.720 ;
        RECT  5.480 2.600 7.000 2.760 ;
        RECT  6.840 0.780 7.000 2.760 ;
        RECT  5.480 0.760 5.640 2.760 ;
        RECT  4.600 0.760 4.760 2.300 ;
        RECT  4.600 0.760 5.640 0.920 ;
        RECT  5.800 0.440 5.960 2.300 ;
        RECT  3.520 0.440 3.680 2.120 ;
        RECT  3.520 0.440 5.960 0.600 ;
        RECT  2.880 2.600 5.320 2.760 ;
        RECT  5.160 1.080 5.320 2.760 ;
        RECT  2.880 0.760 3.040 2.760 ;
        RECT  2.800 0.760 3.040 1.040 ;
        RECT  3.200 2.280 4.240 2.440 ;
        RECT  4.080 0.780 4.240 2.440 ;
        RECT  1.140 2.160 2.300 2.320 ;
        RECT  2.140 0.440 2.300 2.320 ;
        RECT  3.200 0.440 3.360 2.440 ;
        RECT  1.140 0.920 2.300 1.080 ;
        RECT  1.140 0.760 1.420 1.080 ;
        RECT  2.140 0.440 3.360 0.600 ;
        RECT  0.720 2.480 2.720 2.640 ;
        RECT  2.460 2.360 2.720 2.640 ;
        RECT  0.720 0.920 0.880 2.640 ;
    END
END XOR3EHD

MACRO XOR4EHD
    CLASS CORE ;
    FOREIGN XOR4EHD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.000 BY 3.200 ;
    SYMMETRY x y   ;
    SITE core ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  7.700 0.900 7.900 2.750 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  11.300 1.640 11.500 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  10.900 1.240 11.100 1.880 ;
        RECT  10.820 1.240 11.100 1.520 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.500 1.640 0.700 2.280 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.900 1.240 1.180 1.520 ;
        RECT  0.900 1.240 1.100 1.880 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.440 -0.280 3.720 0.400 ;
        RECT  6.890 -0.280 7.170 0.400 ;
        RECT  8.210 -0.280 8.490 0.400 ;
        RECT  10.860 -0.280 11.140 1.080 ;
        RECT  0.000 -0.280 12.000 0.280 ;
        RECT  0.860 -0.280 1.140 1.020 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.400 2.800 3.680 3.480 ;
        RECT  6.880 2.800 7.160 3.480 ;
        RECT  8.210 2.800 8.490 3.480 ;
        RECT  11.040 2.800 11.320 3.480 ;
        RECT  0.000 2.920 12.000 3.480 ;
        RECT  0.680 2.800 0.960 3.480 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  10.080 2.600 10.880 2.760 ;
        RECT  11.720 0.800 11.880 2.640 ;
        RECT  10.720 2.480 11.880 2.640 ;
        RECT  11.660 2.320 11.880 2.640 ;
        RECT  10.080 1.720 10.240 2.760 ;
        RECT  9.020 1.720 9.300 1.940 ;
        RECT  9.020 1.720 10.240 1.880 ;
        RECT  11.660 0.800 11.880 1.080 ;
        RECT  10.400 1.320 10.560 2.440 ;
        RECT  8.720 1.200 8.920 1.520 ;
        RECT  8.720 1.320 10.570 1.480 ;
        RECT  10.120 0.780 10.280 1.480 ;
        RECT  8.760 2.600 9.920 2.760 ;
        RECT  9.760 2.140 9.920 2.760 ;
        RECT  8.060 2.480 8.920 2.640 ;
        RECT  8.060 0.560 8.220 2.640 ;
        RECT  9.360 0.880 9.640 1.040 ;
        RECT  9.360 0.560 9.520 1.040 ;
        RECT  6.450 0.560 9.520 0.720 ;
        RECT  6.450 0.440 6.730 0.720 ;
        RECT  9.100 2.120 9.380 2.360 ;
        RECT  8.380 2.120 9.380 2.280 ;
        RECT  8.380 0.880 8.540 2.280 ;
        RECT  8.380 0.880 9.120 1.040 ;
        RECT  4.480 2.600 6.670 2.760 ;
        RECT  7.380 1.400 7.540 2.640 ;
        RECT  6.510 2.480 7.540 2.640 ;
        RECT  5.410 2.100 5.570 2.760 ;
        RECT  4.480 0.920 4.640 2.760 ;
        RECT  4.480 0.920 4.890 1.080 ;
        RECT  4.730 0.440 4.890 1.080 ;
        RECT  5.430 0.880 5.970 1.040 ;
        RECT  5.430 0.440 5.590 1.040 ;
        RECT  4.730 0.440 5.590 0.600 ;
        RECT  5.950 2.120 6.230 2.320 ;
        RECT  5.950 2.120 7.080 2.280 ;
        RECT  6.920 0.880 7.080 2.280 ;
        RECT  6.210 0.880 7.080 1.040 ;
        RECT  4.800 1.320 4.960 2.380 ;
        RECT  6.570 1.320 6.730 1.800 ;
        RECT  4.800 1.320 6.730 1.480 ;
        RECT  5.050 0.780 5.210 1.480 ;
        RECT  5.170 1.760 6.310 1.920 ;
        RECT  4.130 0.580 4.290 2.230 ;
        RECT  4.130 1.480 4.320 1.760 ;
        RECT  2.080 2.600 3.240 2.760 ;
        RECT  3.810 0.560 3.970 2.640 ;
        RECT  3.080 2.480 3.970 2.640 ;
        RECT  2.080 2.140 2.240 2.760 ;
        RECT  2.360 0.880 2.640 1.040 ;
        RECT  2.480 0.560 2.640 1.040 ;
        RECT  2.480 0.560 3.970 0.720 ;
        RECT  2.620 2.120 2.900 2.360 ;
        RECT  2.620 2.120 3.600 2.280 ;
        RECT  3.440 0.880 3.600 2.280 ;
        RECT  2.880 0.880 3.600 1.040 ;
        RECT  1.440 1.320 1.600 2.420 ;
        RECT  3.020 1.200 3.280 1.520 ;
        RECT  1.430 1.320 3.280 1.480 ;
        RECT  1.660 0.900 1.940 1.480 ;
        RECT  1.120 2.600 1.920 2.760 ;
        RECT  1.760 1.720 1.920 2.760 ;
        RECT  0.120 2.480 1.280 2.640 ;
        RECT  0.120 2.320 0.340 2.640 ;
        RECT  0.120 0.800 0.280 2.640 ;
        RECT  2.700 1.720 2.980 1.940 ;
        RECT  1.760 1.720 2.980 1.880 ;
        RECT  0.120 0.800 0.340 1.080 ;
    END
END XOR4EHD

END LIBRARY
